
module inside_ ( g_input, e_input, o );
  input [72:0] g_input;
  input [24:0] e_input;
  output o;
  wire   \MULT3/B__[0] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n156, n157, n158, n159, n160, n161, n162, n163, n164,
         n165, n166, n167, n168, n169, n170, n171, n172, n173, n174, n175,
         n176, n177, n178, n179, n180, n181, n182, n183, n184, n185, n186,
         n187, n188, n189, n190, n191, n192, n193, n194, n195, n196, n197,
         n198, n199, n200, n201, n202, n203, n204, n205, n206, n207, n208,
         n209, n210, n211, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234, n235, n236, n237, n238, n239, n240, n241,
         n242, n243, n244, n245, n246, n247, n248, n249, n250, n251, n252,
         n253, n254, n255, n256, n257, n258, n259, n260, n261, n262, n263,
         n264, n265, n266, n267, n268, n269, n270, n271, n272, n273, n274,
         n275, n276, n277, n278, n279, n280, n281, n282, n283, n284, n285,
         n286, n287, n288, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328, n329,
         n330, n331, n332, n333, n334, n335, n336, n337, n338, n339, n340,
         n341, n342, n343, n344, n345, n346, n347, n348, n349, n350, n351,
         n352, n353, n354, n355, n356, n357, n358, n359, n360, n361, n362,
         n363, n364, n365, n366, n367, n368, n369, n370, n371, n372, n373,
         n374, n375, n376, n377, n378, n379, n380, n381, n382, n383, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, n398, n399, n400, n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682, n683, n684, n685, n686, n687, n688, n689, n690, n691, n692,
         n693, n694, n695, n696, n697, n698, n699, n700, n701, n702, n703,
         n704, n705, n706, n707, n708, n709, n710, n711, n712, n713, n714,
         n715, n716, n717, n718, n719, n720, n721, n722, n723, n724, n725,
         n726, n727, n728, n729, n730, n731, n732, n733, n734, n735, n736,
         n737, n738, n739, n740, n741, n742, n743, n744, n745, n746, n747,
         n748, n749, n750, n751, n752, n753, n754, n755, n756, n757, n758,
         n759, n760, n761, n762, n763, n764, n765, n766, n767, n768, n769,
         n770, n771, n772, n773, n774, n775, n776, n777, n778, n779, n780,
         n781, n782, n783, n784, n785, n786, n787, n788, n789, n790, n791,
         n792, n793, n794, n795, n796, n797, n798, n799, n800, n801, n802,
         n803, n804, n805, n806, n807, n808, n809, n810, n811, n812, n813,
         n814, n815, n816, n817, n818, n819, n820, n821, n822, n823, n824,
         n825, n826, n827, n828, n829, n830, n831, n832, n833, n834, n835,
         n836, n837, n838, n839, n840, n841, n842, n843, n844, n845, n846,
         n847, n848, n849, n850, n851, n852, n853, n854, n855, n856, n857,
         n858, n859, n860, n861, n862, n863, n864, n865, n866, n867, n868,
         n869, n870, n871, n872, n873, n874, n875, n876, n877, n878, n879,
         n880, n881, n882, n883, n884, n885, n886, n887, n888, n889, n890,
         n891, n892, n893, n894, n895, n896, n897, n898, n899, n900, n901,
         n902, n903, n904, n905, n906, n907, n908, n909, n910, n911, n912,
         n913, n914, n915, n916, n917, n918, n919, n920, n921, n922, n923,
         n924, n925, n926, n927, n928, n929, n930, n931, n932, n933, n934,
         n935, n936, n937, n938, n939, n940, n941, n942, n943, n944, n945,
         n946, n947, n948, n949, n950, n951, n952, n953, n954, n955, n956,
         n957, n958, n959, n960, n961, n962, n963, n964, n965, n966, n967,
         n968, n969, n970, n971, n972, n973, n974, n975, n976, n977, n978,
         n979, n980, n981, n982, n983, n984, n985, n986, n987, n988, n989,
         n990, n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000,
         n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010,
         n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020,
         n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030,
         n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040,
         n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050,
         n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060,
         n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070,
         n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080,
         n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090,
         n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100,
         n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110,
         n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120,
         n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130,
         n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140,
         n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150,
         n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440,
         n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450,
         n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460,
         n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470,
         n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480,
         n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490,
         n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500,
         n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510,
         n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520,
         n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530,
         n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540,
         n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550,
         n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560,
         n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570,
         n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580,
         n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590,
         n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600,
         n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610,
         n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620,
         n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630,
         n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640,
         n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650,
         n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660,
         n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670,
         n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680,
         n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690,
         n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700,
         n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710,
         n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720,
         n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730,
         n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740,
         n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750,
         n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760,
         n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770,
         n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780,
         n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790,
         n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800,
         n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810,
         n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820,
         n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830,
         n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840,
         n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850,
         n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860,
         n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870,
         n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880,
         n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890,
         n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900,
         n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910,
         n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920,
         n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930,
         n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940,
         n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950,
         n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960,
         n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970,
         n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980,
         n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990,
         n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000,
         n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010,
         n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020,
         n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030,
         n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040,
         n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050,
         n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060,
         n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070,
         n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080,
         n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090,
         n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100,
         n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110,
         n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120,
         n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130,
         n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140,
         n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150,
         n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160,
         n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170,
         n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180,
         n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190,
         n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200,
         n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210,
         n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220,
         n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230,
         n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240,
         n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250,
         n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260,
         n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270,
         n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280,
         n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290,
         n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300,
         n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310,
         n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320,
         n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330,
         n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340,
         n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350,
         n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360,
         n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370,
         n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380,
         n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390,
         n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400,
         n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410,
         n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420,
         n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430,
         n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560,
         n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570,
         n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600,
         n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610,
         n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620,
         n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630,
         n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640,
         n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650,
         n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660,
         n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670,
         n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680,
         n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690,
         n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700,
         n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710,
         n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720,
         n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730,
         n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740,
         n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750,
         n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760,
         n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770,
         n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780,
         n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790,
         n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800,
         n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810,
         n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820,
         n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830,
         n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840,
         n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850,
         n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860,
         n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870,
         n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880,
         n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890,
         n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900,
         n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910,
         n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920,
         n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930,
         n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940,
         n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950,
         n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960,
         n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970,
         n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980,
         n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990,
         n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000,
         n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010,
         n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040,
         n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050,
         n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060,
         n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070,
         n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090,
         n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100,
         n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110,
         n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120,
         n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130,
         n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140,
         n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150,
         n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170,
         n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180,
         n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190,
         n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200,
         n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210,
         n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220,
         n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230,
         n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240,
         n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250,
         n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260,
         n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270,
         n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280,
         n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290,
         n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300,
         n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340,
         n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350,
         n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360,
         n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370,
         n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380,
         n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390,
         n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400,
         n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410,
         n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420,
         n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430,
         n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440,
         n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450,
         n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460,
         n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470,
         n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480,
         n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490,
         n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500,
         n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510,
         n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520,
         n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530,
         n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540,
         n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550,
         n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560,
         n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570,
         n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580,
         n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590,
         n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600,
         n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610,
         n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620,
         n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630,
         n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640,
         n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650,
         n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660,
         n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670,
         n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680,
         n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690,
         n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700,
         n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710,
         n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720,
         n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730,
         n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740,
         n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750,
         n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760,
         n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770,
         n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780,
         n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790,
         n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800,
         n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810,
         n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820,
         n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830,
         n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840,
         n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850,
         n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860,
         n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870,
         n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880,
         n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890,
         n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930,
         n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940,
         n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950,
         n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960,
         n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970,
         n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980,
         n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990,
         n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000,
         n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010,
         n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020,
         n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030,
         n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040,
         n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060,
         n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070,
         n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080,
         n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090,
         n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100,
         n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110,
         n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120,
         n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130,
         n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140,
         n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150,
         n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160,
         n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170,
         n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180,
         n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190,
         n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200,
         n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210,
         n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220,
         n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230,
         n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240,
         n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250,
         n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260,
         n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270,
         n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280,
         n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290,
         n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300,
         n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310,
         n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350,
         n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380,
         n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390,
         n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400,
         n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410,
         n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420,
         n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430,
         n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440,
         n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450,
         n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460,
         n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470,
         n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480,
         n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490,
         n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500,
         n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510,
         n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520,
         n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530,
         n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540,
         n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550,
         n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560,
         n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570,
         n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580,
         n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590,
         n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600,
         n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610,
         n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620,
         n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630,
         n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640,
         n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650,
         n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660,
         n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670,
         n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680,
         n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690,
         n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700,
         n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710,
         n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720,
         n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730,
         n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740,
         n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750,
         n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760,
         n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770,
         n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780,
         n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790,
         n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800,
         n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810,
         n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820,
         n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830,
         n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840,
         n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850,
         n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860,
         n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870,
         n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880,
         n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890,
         n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900,
         n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910,
         n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920,
         n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930,
         n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940,
         n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950,
         n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960,
         n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970,
         n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010,
         n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020,
         n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030,
         n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040,
         n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050,
         n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823, n12824,
         n12825, n12826, n12827, n12828, n12829, n12830, n12831, n12832,
         n12833, n12834, n12835, n12836, n12837, n12838, n12839, n12840,
         n12841, n12842, n12843, n12844, n12845, n12846, n12847, n12848,
         n12849, n12850, n12851, n12852, n12853, n12854, n12855, n12856,
         n12857, n12858, n12859, n12860, n12861, n12862, n12863, n12864,
         n12865, n12866, n12867, n12868, n12869, n12870, n12871, n12872,
         n12873, n12874, n12875, n12876, n12877, n12878, n12879, n12880,
         n12881, n12882, n12883, n12884, n12885, n12886, n12887, n12888,
         n12889, n12890, n12891, n12892, n12893, n12894, n12895, n12896,
         n12897, n12898, n12899, n12900, n12901, n12902, n12903, n12904,
         n12905, n12906, n12907, n12908, n12909, n12910, n12911, n12912,
         n12913, n12914, n12915, n12916, n12917, n12918, n12919, n12920,
         n12921, n12922, n12923, n12924, n12925, n12926, n12927, n12928,
         n12929, n12930, n12931, n12932, n12933, n12934, n12935, n12936,
         n12937, n12938, n12939, n12940, n12941, n12942, n12943, n12944,
         n12945, n12946, n12947, n12948, n12949, n12950, n12951, n12952,
         n12953, n12954, n12955, n12956, n12957, n12958, n12959, n12960,
         n12961, n12962, n12963, n12964, n12965, n12966, n12967, n12968,
         n12969, n12970, n12971, n12972, n12973, n12974, n12975, n12976,
         n12977, n12978, n12979, n12980, n12981, n12982, n12983, n12984,
         n12985, n12986, n12987, n12988, n12989, n12990, n12991, n12992,
         n12993, n12994, n12995, n12996, n12997, n12998, n12999, n13000,
         n13001, n13002, n13003, n13004, n13005, n13006, n13007, n13008,
         n13009, n13010, n13011, n13012, n13013, n13014, n13015, n13016,
         n13017, n13018, n13019, n13020, n13021, n13022, n13023, n13024,
         n13025, n13026, n13027, n13028, n13029, n13030, n13031, n13032,
         n13033, n13034, n13035, n13036, n13037, n13038, n13039, n13040,
         n13041, n13042, n13043, n13044, n13045, n13046, n13047, n13048,
         n13049, n13050, n13051, n13052, n13053, n13054, n13055, n13056,
         n13057, n13058, n13059, n13060, n13061, n13062, n13063, n13064,
         n13065, n13066, n13067, n13068, n13069, n13070, n13071, n13072,
         n13073, n13074, n13075, n13076, n13077, n13078, n13079, n13080,
         n13081, n13082, n13083, n13084, n13085, n13086, n13087, n13088,
         n13089, n13090, n13091, n13092, n13093, n13094, n13095, n13096,
         n13097, n13098, n13099, n13100, n13101, n13102, n13103, n13104,
         n13105, n13106, n13107, n13108, n13109, n13110, n13111, n13112,
         n13113, n13114, n13115, n13116, n13117, n13118, n13119, n13120,
         n13121, n13122, n13123, n13124, n13125, n13126, n13127, n13128,
         n13129, n13130, n13131, n13132, n13133, n13134, n13135, n13136,
         n13137, n13138, n13139, n13140, n13141, n13142, n13143, n13144,
         n13145, n13146, n13147, n13148, n13149, n13150, n13151, n13152,
         n13153, n13154, n13155, n13156, n13157, n13158, n13159, n13160,
         n13161, n13162, n13163, n13164, n13165, n13166, n13167, n13168,
         n13169, n13170, n13171, n13172, n13173, n13174, n13175, n13176,
         n13177, n13178, n13179, n13180, n13181, n13182, n13183, n13184,
         n13185, n13186, n13187, n13188, n13189, n13190, n13191, n13192,
         n13193, n13194, n13195, n13196, n13197, n13198, n13199, n13200,
         n13201, n13202, n13203, n13204, n13205, n13206, n13207, n13208,
         n13209, n13210, n13211, n13212, n13213, n13214, n13215, n13216,
         n13217, n13218, n13219, n13220, n13221, n13222, n13223, n13224,
         n13225, n13226, n13227, n13228, n13229, n13230, n13231, n13232,
         n13233, n13234, n13235, n13236, n13237, n13238, n13239, n13240,
         n13241, n13242, n13243, n13244, n13245, n13246, n13247, n13248,
         n13249, n13250, n13251, n13252, n13253, n13254, n13255, n13256,
         n13257, n13258, n13259, n13260, n13261, n13262, n13263, n13264,
         n13265, n13266, n13267, n13268, n13269, n13270, n13271, n13272,
         n13273, n13274, n13275, n13276, n13277, n13278, n13279, n13280,
         n13281, n13282, n13283, n13284, n13285, n13286, n13287, n13288,
         n13289, n13290, n13291, n13292, n13293, n13294, n13295, n13296,
         n13297, n13298, n13299, n13300, n13301, n13302, n13303, n13304,
         n13305, n13306, n13307, n13308, n13309, n13310, n13311, n13312,
         n13313, n13314, n13315, n13316, n13317, n13318, n13319, n13320,
         n13321, n13322, n13323, n13324, n13325, n13326, n13327, n13328,
         n13329, n13330, n13331, n13332, n13333, n13334, n13335, n13336,
         n13337, n13338, n13339, n13340, n13341, n13342, n13343, n13344,
         n13345, n13346, n13347, n13348, n13349, n13350, n13351, n13352,
         n13353, n13354, n13355, n13356, n13357, n13358, n13359, n13360,
         n13361, n13362, n13363, n13364, n13365, n13366, n13367, n13368,
         n13369, n13370, n13371, n13372, n13373, n13374, n13375, n13376,
         n13377, n13378, n13379, n13380, n13381, n13382, n13383, n13384,
         n13385, n13386, n13387, n13388, n13389, n13390, n13391, n13392,
         n13393, n13394, n13395, n13396, n13397, n13398, n13399, n13400,
         n13401, n13402, n13403, n13404, n13405, n13406, n13407, n13408,
         n13409, n13410, n13411, n13412, n13413, n13414, n13415, n13416,
         n13417, n13418, n13419, n13420, n13421, n13422, n13423, n13424,
         n13425, n13426, n13427, n13428, n13429, n13430, n13431, n13432,
         n13433, n13434, n13435, n13436, n13437, n13438, n13439, n13440,
         n13441, n13442, n13443, n13444, n13445, n13446, n13447, n13448,
         n13449, n13450, n13451, n13452, n13453, n13454, n13455, n13456,
         n13457, n13458, n13459, n13460, n13461, n13462, n13463, n13464,
         n13465, n13466, n13467, n13468, n13469, n13470, n13471, n13472,
         n13473, n13474, n13475, n13476, n13477, n13478, n13479, n13480,
         n13481, n13482, n13483, n13484, n13485, n13486, n13487, n13488,
         n13489, n13490, n13491, n13492, n13493, n13494, n13495, n13496,
         n13497, n13498, n13499, n13500, n13501, n13502, n13503, n13504,
         n13505, n13506, n13507, n13508, n13509, n13510, n13511, n13512,
         n13513, n13514, n13515, n13516, n13517, n13518, n13519, n13520,
         n13521, n13522, n13523, n13524, n13525, n13526, n13527, n13528,
         n13529, n13530, n13531, n13532, n13533, n13534, n13535, n13536,
         n13537, n13538, n13539, n13540, n13541, n13542, n13543, n13544,
         n13545, n13546, n13547, n13548, n13549, n13550, n13551, n13552,
         n13553, n13554, n13555, n13556, n13557, n13558, n13559, n13560,
         n13561, n13562, n13563, n13564, n13565, n13566, n13567, n13568,
         n13569, n13570, n13571, n13572, n13573, n13574, n13575, n13576,
         n13577, n13578, n13579, n13580, n13581, n13582, n13583, n13584,
         n13585, n13586, n13587, n13588, n13589, n13590, n13591, n13592,
         n13593, n13594, n13595, n13596, n13597, n13598, n13599, n13600,
         n13601, n13602, n13603, n13604, n13605, n13606, n13607, n13608,
         n13609, n13610, n13611, n13612, n13613, n13614, n13615, n13616,
         n13617, n13618, n13619, n13620, n13621, n13622, n13623, n13624,
         n13625, n13626, n13627, n13628, n13629, n13630, n13631, n13632,
         n13633, n13634, n13635, n13636, n13637, n13638, n13639, n13640,
         n13641, n13642, n13643, n13644, n13645, n13646, n13647, n13648,
         n13649, n13650, n13651, n13652, n13653, n13654, n13655, n13656,
         n13657, n13658, n13659, n13660, n13661, n13662, n13663, n13664,
         n13665, n13666, n13667, n13668, n13669, n13670, n13671, n13672,
         n13673, n13674, n13675, n13676, n13677, n13678, n13679, n13680,
         n13681, n13682, n13683, n13684, n13685, n13686, n13687, n13688,
         n13689, n13690, n13691, n13692, n13693, n13694, n13695, n13696,
         n13697, n13698, n13699, n13700, n13701, n13702, n13703, n13704,
         n13705, n13706, n13707, n13708, n13709, n13710, n13711, n13712,
         n13713, n13714, n13715, n13716, n13717, n13718, n13719, n13720,
         n13721, n13722, n13723, n13724, n13725, n13726, n13727, n13728,
         n13729, n13730, n13731, n13732, n13733, n13734, n13735, n13736,
         n13737, n13738, n13739, n13740, n13741, n13742, n13743, n13744,
         n13745, n13746, n13747, n13748, n13749, n13750, n13751, n13752,
         n13753, n13754, n13755, n13756, n13757, n13758, n13759, n13760,
         n13761, n13762, n13763, n13764, n13765, n13766, n13767, n13768,
         n13769, n13770, n13771, n13772, n13773, n13774, n13775, n13776,
         n13777, n13778, n13779, n13780, n13781, n13782, n13783, n13784,
         n13785, n13786, n13787, n13788, n13789, n13790, n13791, n13792,
         n13793, n13794, n13795, n13796, n13797, n13798, n13799, n13800,
         n13801, n13802, n13803, n13804, n13805, n13806, n13807, n13808,
         n13809, n13810, n13811, n13812, n13813, n13814, n13815, n13816,
         n13817, n13818, n13819, n13820, n13821, n13822, n13823, n13824,
         n13825, n13826, n13827, n13828, n13829, n13830, n13831, n13832,
         n13833, n13834, n13835, n13836, n13837, n13838, n13839, n13840,
         n13841, n13842, n13843, n13844, n13845, n13846, n13847, n13848,
         n13849, n13850, n13851, n13852, n13853, n13854, n13855, n13856,
         n13857, n13858, n13859, n13860, n13861, n13862, n13863, n13864,
         n13865, n13866, n13867, n13868, n13869, n13870, n13871, n13872,
         n13873, n13874, n13875, n13876, n13877, n13878, n13879, n13880,
         n13881, n13882, n13883, n13884, n13885, n13886, n13887, n13888,
         n13889, n13890, n13891, n13892, n13893, n13894, n13895, n13896,
         n13897, n13898, n13899, n13900, n13901, n13902, n13903, n13904,
         n13905, n13906, n13907, n13908, n13909, n13910, n13911, n13912,
         n13913, n13914, n13915, n13916, n13917, n13918, n13919, n13920,
         n13921, n13922, n13923, n13924, n13925, n13926, n13927, n13928,
         n13929, n13930, n13931, n13932, n13933, n13934, n13935, n13936,
         n13937, n13938, n13939, n13940, n13941, n13942, n13943, n13944,
         n13945, n13946, n13947, n13948, n13949, n13950, n13951, n13952,
         n13953, n13954, n13955, n13956, n13957, n13958, n13959, n13960,
         n13961, n13962, n13963, n13964, n13965, n13966, n13967, n13968,
         n13969, n13970, n13971, n13972, n13973, n13974, n13975, n13976,
         n13977, n13978, n13979, n13980, n13981, n13982, n13983, n13984,
         n13985, n13986, n13987, n13988, n13989, n13990, n13991, n13992,
         n13993, n13994, n13995, n13996, n13997, n13998, n13999, n14000,
         n14001, n14002, n14003, n14004, n14005, n14006, n14007, n14008,
         n14009, n14010, n14011, n14012, n14013, n14014, n14015, n14016,
         n14017, n14018, n14019, n14020, n14021, n14022, n14023, n14024,
         n14025, n14026, n14027, n14028, n14029, n14030, n14031, n14032,
         n14033, n14034, n14035, n14036, n14037, n14038, n14039, n14040,
         n14041, n14042, n14043, n14044, n14045, n14046, n14047, n14048,
         n14049, n14050, n14051, n14052, n14053, n14054, n14055, n14056,
         n14057, n14058, n14059, n14060, n14061, n14062, n14063, n14064,
         n14065, n14066, n14067, n14068, n14069, n14070, n14071, n14072,
         n14073, n14074, n14075, n14076, n14077, n14078, n14079, n14080,
         n14081, n14082, n14083, n14084, n14085, n14086, n14087, n14088,
         n14089, n14090, n14091, n14092, n14093, n14094, n14095, n14096,
         n14097, n14098, n14099, n14100, n14101, n14102, n14103, n14104,
         n14105, n14106, n14107, n14108, n14109, n14110, n14111, n14112,
         n14113, n14114, n14115, n14116, n14117, n14118, n14119, n14120,
         n14121, n14122, n14123, n14124, n14125, n14126, n14127, n14128,
         n14129, n14130, n14131, n14132, n14133, n14134, n14135, n14136,
         n14137, n14138, n14139, n14140, n14141, n14142, n14143, n14144,
         n14145, n14146, n14147, n14148, n14149, n14150, n14151, n14152,
         n14153, n14154, n14155, n14156, n14157, n14158, n14159, n14160,
         n14161, n14162, n14163, n14164, n14165, n14166, n14167, n14168,
         n14169, n14170, n14171, n14172, n14173, n14174, n14175, n14176,
         n14177, n14178, n14179, n14180, n14181, n14182, n14183, n14184,
         n14185, n14186, n14187, n14188, n14189, n14190, n14191, n14192,
         n14193, n14194, n14195, n14196, n14197, n14198, n14199, n14200,
         n14201, n14202, n14203, n14204, n14205, n14206, n14207, n14208,
         n14209, n14210, n14211, n14212, n14213, n14214, n14215, n14216,
         n14217, n14218, n14219, n14220, n14221, n14222, n14223, n14224,
         n14225, n14226, n14227, n14228, n14229, n14230, n14231, n14232,
         n14233, n14234, n14235, n14236, n14237, n14238, n14239, n14240,
         n14241, n14242, n14243, n14244, n14245, n14246, n14247, n14248,
         n14249, n14250, n14251, n14252, n14253, n14254, n14255, n14256,
         n14257, n14258, n14259, n14260, n14261, n14262, n14263, n14264,
         n14265, n14266, n14267, n14268, n14269, n14270, n14271, n14272,
         n14273, n14274, n14275, n14276, n14277, n14278, n14279, n14280,
         n14281, n14282, n14283, n14284, n14285, n14286, n14287, n14288,
         n14289, n14290, n14291, n14292, n14293, n14294, n14295, n14296,
         n14297, n14298, n14299, n14300, n14301, n14302, n14303, n14304,
         n14305, n14306, n14307, n14308, n14309, n14310, n14311, n14312,
         n14313, n14314, n14315, n14316, n14317, n14318, n14319, n14320,
         n14321, n14322, n14323, n14324, n14325, n14326, n14327, n14328,
         n14329, n14330, n14331, n14332, n14333, n14334, n14335, n14336,
         n14337, n14338, n14339, n14340, n14341, n14342, n14343, n14344,
         n14345, n14346, n14347, n14348, n14349, n14350, n14351, n14352,
         n14353, n14354, n14355, n14356, n14357, n14358, n14359, n14360,
         n14361, n14362, n14363, n14364, n14365, n14366, n14367, n14368,
         n14369, n14370, n14371, n14372, n14373, n14374, n14375, n14376,
         n14377, n14378, n14379, n14380, n14381, n14382, n14383, n14384,
         n14385, n14386, n14387, n14388, n14389, n14390, n14391, n14392,
         n14393, n14394, n14395, n14396, n14397, n14398, n14399, n14400,
         n14401, n14402, n14403, n14404, n14405, n14406, n14407, n14408,
         n14409, n14410, n14411, n14412, n14413, n14414, n14415, n14416,
         n14417, n14418, n14419, n14420, n14421, n14422, n14423, n14424,
         n14425, n14426, n14427, n14428, n14429, n14430, n14431, n14432,
         n14433, n14434, n14435, n14436, n14437, n14438, n14439, n14440,
         n14441, n14442, n14443, n14444, n14445, n14446, n14447, n14448,
         n14449, n14450, n14451, n14452, n14453, n14454, n14455, n14456,
         n14457, n14458, n14459, n14460, n14461, n14462, n14463, n14464,
         n14465, n14466, n14467, n14468, n14469, n14470, n14471, n14472,
         n14473, n14474, n14475, n14476, n14477, n14478, n14479, n14480,
         n14481, n14482, n14483, n14484, n14485, n14486, n14487, n14488,
         n14489, n14490, n14491, n14492, n14493, n14494, n14495, n14496,
         n14497, n14498, n14499, n14500, n14501, n14502, n14503, n14504,
         n14505, n14506, n14507, n14508, n14509, n14510, n14511, n14512,
         n14513, n14514, n14515, n14516, n14517, n14518, n14519, n14520,
         n14521, n14522, n14523, n14524, n14525, n14526, n14527, n14528,
         n14529, n14530, n14531, n14532, n14533, n14534, n14535, n14536,
         n14537, n14538, n14539, n14540, n14541, n14542, n14543, n14544,
         n14545, n14546, n14547, n14548, n14549, n14550, n14551, n14552,
         n14553, n14554, n14555, n14556, n14557, n14558, n14559, n14560,
         n14561, n14562, n14563, n14564, n14565, n14566, n14567, n14568,
         n14569, n14570, n14571, n14572, n14573, n14574, n14575, n14576,
         n14577, n14578, n14579, n14580, n14581, n14582, n14583, n14584,
         n14585, n14586, n14587, n14588, n14589, n14590, n14591, n14592,
         n14593, n14594, n14595, n14596, n14597, n14598, n14599, n14600,
         n14601, n14602, n14603, n14604, n14605, n14606, n14607, n14608,
         n14609, n14610, n14611, n14612, n14613, n14614, n14615, n14616,
         n14617, n14618, n14619, n14620, n14621, n14622, n14623, n14624,
         n14625, n14626, n14627, n14628, n14629, n14630, n14631, n14632,
         n14633, n14634, n14635, n14636, n14637, n14638, n14639, n14640,
         n14641, n14642, n14643, n14644, n14645, n14646, n14647, n14648,
         n14649, n14650, n14651, n14652, n14653, n14654, n14655, n14656,
         n14657, n14658, n14659, n14660, n14661, n14662, n14663, n14664,
         n14665, n14666, n14667, n14668, n14669, n14670, n14671, n14672,
         n14673, n14674, n14675, n14676, n14677, n14678, n14679, n14680,
         n14681, n14682, n14683, n14684, n14685, n14686, n14687, n14688,
         n14689, n14690, n14691, n14692, n14693, n14694, n14695, n14696,
         n14697, n14698, n14699, n14700, n14701, n14702, n14703, n14704,
         n14705, n14706, n14707, n14708, n14709, n14710, n14711, n14712,
         n14713, n14714, n14715, n14716, n14717, n14718, n14719, n14720,
         n14721, n14722, n14723, n14724, n14725, n14726, n14727, n14728,
         n14729, n14730, n14731, n14732, n14733, n14734, n14735, n14736,
         n14737, n14738, n14739, n14740, n14741, n14742, n14743, n14744,
         n14745, n14746, n14747, n14748, n14749, n14750, n14751, n14752,
         n14753, n14754, n14755, n14756, n14757, n14758, n14759, n14760,
         n14761, n14762, n14763, n14764, n14765, n14766, n14767, n14768,
         n14769, n14770, n14771, n14772, n14773, n14774, n14775, n14776,
         n14777, n14778, n14779, n14780, n14781, n14782, n14783, n14784,
         n14785, n14786, n14787, n14788, n14789, n14790, n14791, n14792,
         n14793, n14794, n14795, n14796, n14797, n14798, n14799, n14800,
         n14801, n14802, n14803, n14804, n14805, n14806, n14807, n14808,
         n14809, n14810, n14811, n14812, n14813, n14814, n14815, n14816,
         n14817, n14818, n14819, n14820, n14821, n14822, n14823, n14824,
         n14825, n14826, n14827, n14828, n14829, n14830, n14831, n14832,
         n14833, n14834, n14835, n14836, n14837, n14838, n14839, n14840,
         n14841, n14842, n14843, n14844, n14845, n14846, n14847, n14848,
         n14849, n14850, n14851, n14852, n14853, n14854, n14855, n14856,
         n14857, n14858, n14859, n14860, n14861, n14862, n14863, n14864,
         n14865, n14866, n14867, n14868, n14869, n14870, n14871, n14872,
         n14873, n14874, n14875, n14876, n14877, n14878, n14879, n14880,
         n14881, n14882, n14883, n14884, n14885, n14886, n14887, n14888,
         n14889, n14890, n14891, n14892, n14893, n14894, n14895, n14896,
         n14897, n14898, n14899, n14900, n14901, n14902, n14903, n14904,
         n14905, n14906, n14907, n14908, n14909, n14910, n14911, n14912,
         n14913, n14914, n14915, n14916, n14917, n14918, n14919, n14920,
         n14921, n14922, n14923, n14924, n14925, n14926, n14927, n14928,
         n14929, n14930, n14931, n14932, n14933, n14934, n14935, n14936,
         n14937, n14938, n14939, n14940, n14941, n14942, n14943, n14944,
         n14945, n14946, n14947, n14948, n14949, n14950, n14951, n14952,
         n14953, n14954, n14955, n14956, n14957, n14958, n14959, n14960,
         n14961, n14962, n14963, n14964, n14965, n14966, n14967, n14968,
         n14969, n14970, n14971, n14972, n14973, n14974, n14975, n14976,
         n14977, n14978, n14979, n14980, n14981, n14982, n14983, n14984,
         n14985, n14986, n14987, n14988, n14989, n14990, n14991, n14992,
         n14993, n14994, n14995, n14996, n14997, n14998, n14999, n15000,
         n15001, n15002, n15003, n15004, n15005, n15006, n15007, n15008,
         n15009, n15010, n15011, n15012, n15013, n15014, n15015, n15016,
         n15017, n15018, n15019, n15020, n15021, n15022, n15023, n15024,
         n15025, n15026, n15027, n15028, n15029, n15030, n15031, n15032,
         n15033, n15034, n15035, n15036, n15037, n15038, n15039, n15040,
         n15041, n15042, n15043, n15044, n15045, n15046, n15047, n15048,
         n15049, n15050, n15051, n15052, n15053, n15054, n15055, n15056,
         n15057, n15058, n15059, n15060, n15061, n15062, n15063, n15064,
         n15065, n15066, n15067, n15068, n15069, n15070, n15071, n15072,
         n15073, n15074, n15075, n15076, n15077, n15078, n15079, n15080,
         n15081, n15082, n15083, n15084, n15085, n15086, n15087, n15088,
         n15089, n15090, n15091, n15092, n15093, n15094, n15095, n15096,
         n15097, n15098, n15099, n15100, n15101, n15102, n15103, n15104,
         n15105, n15106, n15107, n15108, n15109, n15110, n15111, n15112,
         n15113, n15114, n15115, n15116, n15117, n15118, n15119, n15120,
         n15121, n15122, n15123, n15124, n15125, n15126, n15127, n15128,
         n15129, n15130, n15131, n15132, n15133, n15134, n15135, n15136,
         n15137, n15138, n15139, n15140, n15141, n15142, n15143, n15144,
         n15145, n15146, n15147, n15148, n15149, n15150, n15151, n15152,
         n15153, n15154, n15155, n15156, n15157, n15158, n15159, n15160,
         n15161, n15162, n15163, n15164, n15165, n15166, n15167, n15168,
         n15169, n15170, n15171, n15172, n15173, n15174, n15175, n15176,
         n15177, n15178, n15179, n15180, n15181, n15182, n15183, n15184,
         n15185, n15186, n15187, n15188, n15189, n15190, n15191, n15192,
         n15193, n15194, n15195, n15196, n15197, n15198, n15199, n15200,
         n15201, n15202, n15203, n15204, n15205, n15206, n15207, n15208,
         n15209, n15210, n15211, n15212, n15213, n15214, n15215, n15216,
         n15217, n15218, n15219, n15220, n15221, n15222, n15223, n15224,
         n15225, n15226, n15227, n15228, n15229, n15230, n15231, n15232,
         n15233, n15234, n15235, n15236, n15237, n15238, n15239, n15240,
         n15241, n15242, n15243, n15244, n15245, n15246, n15247, n15248,
         n15249, n15250, n15251, n15252, n15253, n15254, n15255, n15256,
         n15257, n15258, n15259, n15260, n15261, n15262, n15263, n15264,
         n15265, n15266, n15267, n15268, n15269, n15270, n15271, n15272,
         n15273, n15274, n15275, n15276, n15277, n15278, n15279, n15280,
         n15281, n15282, n15283, n15284, n15285, n15286, n15287, n15288,
         n15289, n15290, n15291, n15292, n15293, n15294, n15295, n15296,
         n15297, n15298, n15299, n15300, n15301, n15302, n15303, n15304,
         n15305, n15306, n15307, n15308, n15309, n15310, n15311, n15312,
         n15313, n15314, n15315, n15316, n15317, n15318, n15319, n15320,
         n15321, n15322, n15323, n15324, n15325, n15326, n15327, n15328,
         n15329, n15330, n15331, n15332, n15333, n15334, n15335, n15336,
         n15337, n15338, n15339, n15340, n15341, n15342, n15343, n15344,
         n15345, n15346, n15347, n15348, n15349, n15350, n15351, n15352,
         n15353, n15354, n15355, n15356, n15357, n15358, n15359, n15360,
         n15361, n15362, n15363, n15364, n15365, n15366, n15367, n15368,
         n15369, n15370, n15371, n15372, n15373, n15374, n15375, n15376,
         n15377, n15378, n15379, n15380, n15381, n15382, n15383, n15384,
         n15385, n15386, n15387, n15388, n15389, n15390, n15391, n15392,
         n15393, n15394, n15395, n15396, n15397, n15398, n15399, n15400,
         n15401, n15402, n15403, n15404, n15405, n15406, n15407, n15408,
         n15409, n15410, n15411, n15412, n15413, n15414, n15415, n15416,
         n15417, n15418, n15419, n15420, n15421, n15422, n15423, n15424,
         n15425, n15426, n15427, n15428, n15429, n15430, n15431, n15432,
         n15433, n15434, n15435, n15436, n15437, n15438, n15439, n15440,
         n15441, n15442, n15443, n15444, n15445, n15446, n15447, n15448,
         n15449, n15450, n15451, n15452, n15453, n15454, n15455, n15456,
         n15457, n15458, n15459, n15460, n15461, n15462, n15463, n15464,
         n15465, n15466, n15467, n15468, n15469, n15470, n15471, n15472,
         n15473, n15474, n15475, n15476, n15477, n15478, n15479, n15480,
         n15481, n15482, n15483, n15484, n15485, n15486, n15487, n15488,
         n15489, n15490, n15491, n15492, n15493, n15494, n15495, n15496,
         n15497, n15498, n15499, n15500, n15501, n15502, n15503, n15504,
         n15505, n15506, n15507, n15508, n15509, n15510, n15511, n15512,
         n15513, n15514, n15515, n15516, n15517, n15518, n15519, n15520,
         n15521, n15522, n15523, n15524, n15525, n15526, n15527, n15528,
         n15529, n15530, n15531, n15532, n15533, n15534, n15535, n15536,
         n15537, n15538, n15539, n15540, n15541, n15542, n15543, n15544,
         n15545, n15546, n15547, n15548, n15549, n15550, n15551, n15552,
         n15553, n15554, n15555, n15556, n15557, n15558, n15559, n15560,
         n15561, n15562, n15563, n15564, n15565, n15566, n15567, n15568,
         n15569, n15570, n15571, n15572, n15573, n15574, n15575, n15576,
         n15577, n15578, n15579, n15580, n15581, n15582, n15583, n15584,
         n15585, n15586, n15587, n15588, n15589, n15590, n15591, n15592,
         n15593, n15594, n15595, n15596, n15597, n15598, n15599, n15600,
         n15601, n15602, n15603, n15604, n15605, n15606, n15607, n15608,
         n15609, n15610, n15611, n15612, n15613, n15614, n15615, n15616,
         n15617, n15618, n15619, n15620, n15621, n15622, n15623, n15624,
         n15625, n15626, n15627, n15628, n15629, n15630, n15631, n15632,
         n15633, n15634, n15635, n15636, n15637, n15638, n15639, n15640,
         n15641, n15642, n15643, n15644, n15645, n15646, n15647, n15648,
         n15649, n15650, n15651, n15652, n15653, n15654, n15655, n15656,
         n15657, n15658, n15659, n15660, n15661, n15662, n15663, n15664,
         n15665, n15666, n15667, n15668, n15669, n15670, n15671, n15672,
         n15673, n15674, n15675, n15676, n15677, n15678, n15679, n15680,
         n15681, n15682, n15683, n15684, n15685, n15686, n15687, n15688,
         n15689, n15690, n15691, n15692, n15693, n15694, n15695, n15696,
         n15697, n15698, n15699, n15700, n15701, n15702, n15703, n15704,
         n15705, n15706, n15707, n15708, n15709, n15710, n15711, n15712,
         n15713, n15714, n15715, n15716, n15717, n15718, n15719, n15720,
         n15721, n15722, n15723, n15724, n15725, n15726, n15727, n15728,
         n15729, n15730, n15731, n15732, n15733, n15734, n15735, n15736,
         n15737, n15738, n15739, n15740, n15741, n15742, n15743, n15744,
         n15745, n15746, n15747, n15748, n15749, n15750, n15751, n15752,
         n15753, n15754, n15755, n15756, n15757, n15758, n15759, n15760,
         n15761, n15762, n15763, n15764, n15765, n15766, n15767, n15768,
         n15769, n15770, n15771, n15772, n15773, n15774, n15775, n15776,
         n15777, n15778, n15779, n15780, n15781, n15782, n15783, n15784,
         n15785, n15786, n15787, n15788, n15789, n15790, n15791, n15792,
         n15793, n15794, n15795, n15796, n15797, n15798, n15799, n15800,
         n15801, n15802, n15803, n15804, n15805, n15806, n15807, n15808,
         n15809, n15810, n15811, n15812, n15813, n15814, n15815, n15816,
         n15817, n15818, n15819, n15820, n15821, n15822, n15823, n15824,
         n15825, n15826, n15827, n15828, n15829, n15830, n15831, n15832,
         n15833, n15834, n15835, n15836, n15837, n15838, n15839, n15840,
         n15841, n15842, n15843, n15844, n15845, n15846, n15847, n15848,
         n15849, n15850, n15851, n15852, n15853, n15854, n15855, n15856,
         n15857, n15858, n15859, n15860, n15861, n15862, n15863, n15864,
         n15865, n15866, n15867, n15868, n15869, n15870, n15871, n15872,
         n15873, n15874, n15875, n15876, n15877, n15878, n15879, n15880,
         n15881, n15882, n15883, n15884, n15885, n15886, n15887, n15888,
         n15889, n15890, n15891, n15892, n15893, n15894, n15895, n15896,
         n15897, n15898, n15899, n15900, n15901, n15902, n15903, n15904,
         n15905, n15906, n15907, n15908, n15909, n15910, n15911, n15912,
         n15913, n15914, n15915, n15916, n15917, n15918, n15919, n15920,
         n15921, n15922, n15923, n15924, n15925, n15926, n15927, n15928,
         n15929, n15930, n15931, n15932, n15933, n15934, n15935, n15936,
         n15937, n15938, n15939, n15940, n15941, n15942, n15943, n15944,
         n15945, n15946, n15947, n15948, n15949, n15950, n15951, n15952,
         n15953, n15954, n15955, n15956, n15957, n15958, n15959, n15960,
         n15961, n15962, n15963, n15964, n15965, n15966, n15967, n15968,
         n15969, n15970, n15971, n15972, n15973, n15974, n15975, n15976,
         n15977, n15978, n15979, n15980, n15981, n15982, n15983, n15984,
         n15985, n15986, n15987, n15988, n15989, n15990, n15991, n15992,
         n15993, n15994, n15995, n15996, n15997, n15998, n15999, n16000,
         n16001, n16002, n16003, n16004, n16005, n16006, n16007, n16008,
         n16009, n16010, n16011, n16012, n16013, n16014, n16015, n16016,
         n16017, n16018, n16019, n16020, n16021, n16022, n16023, n16024,
         n16025, n16026, n16027, n16028, n16029, n16030, n16031, n16032,
         n16033, n16034, n16035, n16036, n16037, n16038, n16039, n16040,
         n16041, n16042, n16043, n16044, n16045, n16046, n16047, n16048,
         n16049, n16050, n16051, n16052, n16053, n16054, n16055, n16056,
         n16057, n16058, n16059, n16060, n16061, n16062, n16063, n16064,
         n16065, n16066, n16067, n16068, n16069, n16070, n16071, n16072,
         n16073, n16074, n16075, n16076, n16077, n16078, n16079, n16080,
         n16081, n16082, n16083, n16084, n16085, n16086, n16087, n16088,
         n16089, n16090, n16091, n16092, n16093, n16094, n16095, n16096,
         n16097, n16098, n16099, n16100, n16101, n16102, n16103, n16104,
         n16105, n16106, n16107, n16108, n16109, n16110, n16111, n16112,
         n16113, n16114, n16115, n16116, n16117, n16118, n16119, n16120,
         n16121, n16122, n16123, n16124, n16125, n16126, n16127, n16128,
         n16129, n16130, n16131, n16132, n16133, n16134, n16135, n16136,
         n16137, n16138, n16139, n16140, n16141, n16142, n16143, n16144,
         n16145, n16146, n16147, n16148, n16149, n16150, n16151, n16152,
         n16153, n16154, n16155, n16156, n16157, n16158, n16159, n16160,
         n16161, n16162, n16163, n16164, n16165, n16166, n16167, n16168,
         n16169, n16170, n16171, n16172, n16173, n16174, n16175, n16176,
         n16177, n16178, n16179, n16180, n16181, n16182, n16183, n16184,
         n16185, n16186, n16187, n16188, n16189, n16190, n16191, n16192,
         n16193, n16194, n16195, n16196, n16197, n16198, n16199, n16200,
         n16201, n16202, n16203, n16204, n16205, n16206, n16207, n16208,
         n16209, n16210, n16211, n16212, n16213, n16214, n16215, n16216,
         n16217, n16218, n16219, n16220, n16221, n16222, n16223, n16224,
         n16225, n16226, n16227, n16228, n16229, n16230, n16231, n16232,
         n16233, n16234, n16235, n16236, n16237, n16238, n16239, n16240,
         n16241, n16242, n16243, n16244, n16245, n16246, n16247, n16248,
         n16249, n16250, n16251, n16252, n16253, n16254, n16255, n16256,
         n16257, n16258, n16259, n16260, n16261, n16262, n16263, n16264,
         n16265, n16266, n16267, n16268, n16269, n16270, n16271, n16272,
         n16273, n16274, n16275, n16276, n16277, n16278, n16279, n16280,
         n16281, n16282, n16283, n16284, n16285, n16286, n16287, n16288,
         n16289, n16290, n16291, n16292, n16293, n16294, n16295, n16296,
         n16297, n16298, n16299, n16300, n16301, n16302, n16303, n16304,
         n16305, n16306, n16307, n16308, n16309, n16310, n16311, n16312,
         n16313, n16314, n16315, n16316, n16317, n16318, n16319, n16320,
         n16321, n16322, n16323, n16324, n16325, n16326, n16327, n16328,
         n16329, n16330, n16331, n16332, n16333, n16334, n16335, n16336,
         n16337, n16338, n16339, n16340, n16341, n16342, n16343, n16344,
         n16345, n16346, n16347, n16348, n16349, n16350, n16351, n16352,
         n16353, n16354, n16355, n16356, n16357, n16358, n16359, n16360,
         n16361, n16362, n16363, n16364, n16365, n16366, n16367, n16368,
         n16369, n16370, n16371, n16372, n16373, n16374, n16375, n16376,
         n16377, n16378, n16379, n16380, n16381, n16382, n16383, n16384,
         n16385, n16386, n16387, n16388, n16389, n16390, n16391, n16392,
         n16393, n16394, n16395, n16396, n16397, n16398, n16399, n16400,
         n16401, n16402, n16403, n16404, n16405, n16406, n16407, n16408,
         n16409, n16410, n16411, n16412, n16413, n16414, n16415, n16416,
         n16417, n16418, n16419, n16420, n16421, n16422, n16423, n16424,
         n16425, n16426, n16427, n16428, n16429, n16430, n16431, n16432,
         n16433, n16434, n16435, n16436, n16437, n16438, n16439, n16440,
         n16441, n16442, n16443, n16444, n16445, n16446, n16447, n16448,
         n16449, n16450, n16451, n16452, n16453, n16454, n16455, n16456,
         n16457, n16458, n16459, n16460, n16461, n16462, n16463, n16464,
         n16465, n16466, n16467, n16468, n16469, n16470, n16471, n16472,
         n16473, n16474, n16475, n16476, n16477, n16478, n16479, n16480,
         n16481, n16482, n16483, n16484, n16485, n16486, n16487, n16488,
         n16489, n16490, n16491, n16492, n16493, n16494, n16495, n16496,
         n16497, n16498, n16499, n16500, n16501, n16502, n16503, n16504,
         n16505, n16506, n16507, n16508, n16509, n16510, n16511, n16512,
         n16513, n16514, n16515, n16516, n16517, n16518, n16519, n16520,
         n16521, n16522, n16523, n16524, n16525, n16526, n16527, n16528,
         n16529, n16530, n16531, n16532, n16533, n16534, n16535, n16536,
         n16537, n16538, n16539, n16540, n16541, n16542, n16543, n16544,
         n16545, n16546, n16547, n16548, n16549, n16550, n16551, n16552,
         n16553, n16554, n16555, n16556, n16557, n16558, n16559, n16560,
         n16561, n16562, n16563, n16564, n16565, n16566, n16567, n16568,
         n16569, n16570, n16571, n16572, n16573, n16574, n16575, n16576,
         n16577, n16578, n16579, n16580, n16581, n16582, n16583, n16584,
         n16585, n16586, n16587, n16588, n16589, n16590, n16591, n16592,
         n16593, n16594, n16595, n16596, n16597, n16598, n16599, n16600,
         n16601, n16602, n16603, n16604, n16605, n16606, n16607, n16608,
         n16609, n16610, n16611, n16612, n16613, n16614, n16615, n16616,
         n16617, n16618, n16619, n16620, n16621, n16622, n16623, n16624,
         n16625, n16626, n16627, n16628, n16629, n16630, n16631, n16632,
         n16633, n16634, n16635, n16636, n16637, n16638, n16639, n16640,
         n16641, n16642, n16643, n16644, n16645, n16646, n16647, n16648,
         n16649, n16650, n16651, n16652, n16653, n16654, n16655, n16656,
         n16657, n16658, n16659, n16660, n16661, n16662, n16663, n16664,
         n16665, n16666, n16667, n16668, n16669, n16670, n16671, n16672,
         n16673, n16674, n16675, n16676, n16677, n16678, n16679, n16680,
         n16681, n16682, n16683, n16684, n16685, n16686, n16687, n16688,
         n16689, n16690, n16691, n16692, n16693, n16694, n16695, n16696,
         n16697, n16698, n16699, n16700, n16701, n16702, n16703, n16704,
         n16705, n16706, n16707, n16708, n16709, n16710, n16711, n16712,
         n16713, n16714, n16715, n16716, n16717, n16718, n16719, n16720,
         n16721, n16722, n16723, n16724, n16725, n16726, n16727, n16728,
         n16729, n16730, n16731, n16732, n16733, n16734, n16735, n16736,
         n16737, n16738, n16739, n16740, n16741, n16742, n16743, n16744,
         n16745, n16746, n16747, n16748, n16749, n16750, n16751, n16752,
         n16753, n16754, n16755, n16756, n16757, n16758, n16759, n16760,
         n16761, n16762, n16763, n16764, n16765, n16766, n16767, n16768,
         n16769, n16770, n16771, n16772, n16773, n16774, n16775, n16776,
         n16777, n16778, n16779, n16780, n16781, n16782, n16783, n16784,
         n16785, n16786, n16787, n16788, n16789, n16790, n16791, n16792,
         n16793, n16794, n16795, n16796, n16797, n16798, n16799, n16800,
         n16801, n16802, n16803, n16804, n16805, n16806, n16807, n16808,
         n16809, n16810, n16811, n16812, n16813, n16814, n16815, n16816,
         n16817, n16818, n16819, n16820, n16821, n16822, n16823, n16824,
         n16825, n16826, n16827, n16828, n16829, n16830, n16831, n16832,
         n16833, n16834, n16835, n16836, n16837, n16838, n16839, n16840,
         n16841, n16842, n16843, n16844, n16845, n16846, n16847, n16848,
         n16849, n16850, n16851, n16852, n16853, n16854, n16855, n16856,
         n16857, n16858, n16859, n16860, n16861, n16862, n16863, n16864,
         n16865, n16866, n16867, n16868, n16869, n16870, n16871, n16872,
         n16873, n16874, n16875, n16876, n16877, n16878, n16879, n16880,
         n16881, n16882, n16883, n16884, n16885, n16886, n16887, n16888,
         n16889, n16890, n16891, n16892, n16893, n16894, n16895, n16896,
         n16897, n16898, n16899, n16900, n16901, n16902, n16903, n16904,
         n16905, n16906, n16907, n16908, n16909, n16910, n16911, n16912,
         n16913, n16914, n16915, n16916, n16917, n16918, n16919, n16920,
         n16921, n16922, n16923, n16924, n16925, n16926, n16927, n16928,
         n16929, n16930, n16931, n16932, n16933, n16934, n16935, n16936,
         n16937, n16938, n16939, n16940, n16941, n16942, n16943, n16944,
         n16945, n16946, n16947, n16948, n16949, n16950, n16951, n16952,
         n16953, n16954, n16955, n16956, n16957, n16958, n16959, n16960,
         n16961, n16962, n16963, n16964, n16965, n16966, n16967, n16968,
         n16969, n16970, n16971, n16972, n16973, n16974, n16975, n16976,
         n16977, n16978, n16979, n16980, n16981, n16982, n16983, n16984,
         n16985, n16986, n16987, n16988, n16989, n16990, n16991, n16992,
         n16993, n16994, n16995, n16996, n16997, n16998, n16999, n17000,
         n17001, n17002, n17003, n17004, n17005, n17006, n17007, n17008,
         n17009, n17010, n17011, n17012, n17013, n17014, n17015, n17016,
         n17017, n17018, n17019, n17020, n17021, n17022, n17023, n17024,
         n17025, n17026, n17027, n17028, n17029, n17030, n17031, n17032,
         n17033, n17034, n17035, n17036, n17037, n17038, n17039, n17040,
         n17041, n17042, n17043, n17044, n17045, n17046, n17047, n17048,
         n17049, n17050, n17051, n17052, n17053, n17054, n17055, n17056,
         n17057, n17058, n17059, n17060, n17061, n17062, n17063, n17064,
         n17065, n17066, n17067, n17068, n17069, n17070, n17071, n17072,
         n17073, n17074, n17075, n17076, n17077, n17078, n17079, n17080,
         n17081, n17082, n17083, n17084, n17085, n17086, n17087, n17088,
         n17089, n17090, n17091, n17092, n17093, n17094, n17095, n17096,
         n17097, n17098, n17099, n17100, n17101, n17102, n17103, n17104,
         n17105, n17106, n17107, n17108, n17109, n17110, n17111, n17112,
         n17113, n17114, n17115, n17116, n17117, n17118, n17119, n17120,
         n17121, n17122, n17123, n17124, n17125, n17126, n17127, n17128,
         n17129, n17130, n17131, n17132, n17133, n17134, n17135, n17136,
         n17137, n17138, n17139, n17140, n17141, n17142, n17143, n17144,
         n17145, n17146, n17147, n17148, n17149, n17150, n17151, n17152,
         n17153, n17154, n17155, n17156, n17157, n17158, n17159, n17160,
         n17161, n17162, n17163, n17164, n17165, n17166, n17167, n17168,
         n17169, n17170, n17171, n17172, n17173, n17174, n17175, n17176,
         n17177, n17178, n17179, n17180, n17181, n17182, n17183, n17184,
         n17185, n17186, n17187, n17188, n17189, n17190, n17191, n17192,
         n17193, n17194, n17195, n17196, n17197, n17198, n17199, n17200,
         n17201, n17202, n17203, n17204, n17205, n17206, n17207, n17208,
         n17209, n17210, n17211, n17212, n17213, n17214, n17215, n17216,
         n17217, n17218, n17219, n17220, n17221, n17222, n17223, n17224,
         n17225, n17226, n17227, n17228, n17229, n17230, n17231, n17232,
         n17233, n17234, n17235, n17236, n17237, n17238, n17239, n17240,
         n17241, n17242, n17243, n17244, n17245, n17246, n17247, n17248,
         n17249, n17250, n17251, n17252, n17253, n17254, n17255, n17256,
         n17257, n17258, n17259, n17260, n17261, n17262, n17263, n17264,
         n17265, n17266, n17267, n17268, n17269, n17270, n17271, n17272,
         n17273, n17274, n17275, n17276, n17277, n17278, n17279, n17280,
         n17281, n17282, n17283, n17284, n17285, n17286, n17287, n17288,
         n17289, n17290, n17291, n17292, n17293, n17294, n17295, n17296,
         n17297, n17298, n17299, n17300, n17301, n17302, n17303, n17304,
         n17305, n17306, n17307, n17308, n17309, n17310, n17311, n17312,
         n17313, n17314, n17315, n17316, n17317, n17318, n17319, n17320,
         n17321, n17322, n17323, n17324, n17325, n17326, n17327, n17328,
         n17329, n17330, n17331, n17332, n17333, n17334, n17335, n17336,
         n17337, n17338, n17339, n17340, n17341, n17342, n17343, n17344,
         n17345, n17346, n17347, n17348, n17349, n17350, n17351, n17352,
         n17353, n17354, n17355, n17356, n17357, n17358, n17359, n17360,
         n17361, n17362, n17363, n17364, n17365, n17366, n17367, n17368,
         n17369, n17370, n17371, n17372, n17373, n17374, n17375, n17376,
         n17377, n17378, n17379, n17380, n17381, n17382, n17383, n17384,
         n17385, n17386, n17387, n17388, n17389, n17390, n17391, n17392,
         n17393, n17394, n17395, n17396, n17397, n17398, n17399, n17400,
         n17401, n17402, n17403, n17404, n17405, n17406, n17407, n17408,
         n17409, n17410, n17411, n17412, n17413, n17414, n17415, n17416,
         n17417, n17418, n17419, n17420, n17421, n17422, n17423, n17424,
         n17425, n17426, n17427, n17428, n17429, n17430, n17431, n17432,
         n17433, n17434, n17435, n17436, n17437, n17438, n17439, n17440,
         n17441, n17442, n17443, n17444, n17445, n17446, n17447, n17448,
         n17449, n17450, n17451, n17452, n17453, n17454, n17455, n17456,
         n17457, n17458, n17459, n17460, n17461, n17462, n17463, n17464,
         n17465, n17466, n17467, n17468, n17469, n17470, n17471, n17472,
         n17473, n17474, n17475, n17476, n17477, n17478, n17479, n17480,
         n17481, n17482, n17483, n17484, n17485, n17486, n17487, n17488,
         n17489, n17490, n17491, n17492, n17493, n17494, n17495, n17496,
         n17497, n17498, n17499, n17500, n17501, n17502, n17503, n17504,
         n17505, n17506, n17507, n17508, n17509, n17510, n17511, n17512,
         n17513, n17514, n17515, n17516, n17517, n17518, n17519, n17520,
         n17521, n17522, n17523, n17524, n17525, n17526, n17527, n17528,
         n17529, n17530, n17531, n17532, n17533, n17534, n17535, n17536,
         n17537, n17538, n17539, n17540, n17541, n17542, n17543, n17544,
         n17545, n17546, n17547, n17548, n17549, n17550, n17551, n17552,
         n17553, n17554, n17555, n17556, n17557, n17558, n17559, n17560,
         n17561, n17562, n17563, n17564, n17565, n17566, n17567, n17568,
         n17569, n17570, n17571, n17572, n17573, n17574, n17575, n17576,
         n17577, n17578, n17579, n17580, n17581, n17582, n17583, n17584,
         n17585, n17586, n17587, n17588, n17589, n17590, n17591, n17592,
         n17593, n17594, n17595, n17596, n17597, n17598, n17599, n17600,
         n17601, n17602, n17603, n17604, n17605, n17606, n17607, n17608,
         n17609, n17610, n17611, n17612, n17613, n17614, n17615, n17616,
         n17617, n17618, n17619, n17620, n17621, n17622, n17623, n17624,
         n17625, n17626, n17627, n17628, n17629, n17630, n17631, n17632,
         n17633, n17634, n17635, n17636, n17637, n17638, n17639, n17640,
         n17641, n17642, n17643, n17644, n17645, n17646, n17647, n17648,
         n17649, n17650, n17651, n17652, n17653, n17654, n17655, n17656,
         n17657, n17658, n17659, n17660, n17661, n17662, n17663, n17664,
         n17665, n17666, n17667, n17668, n17669, n17670, n17671, n17672,
         n17673, n17674, n17675, n17676, n17677, n17678, n17679, n17680,
         n17681, n17682, n17683, n17684, n17685, n17686, n17687, n17688,
         n17689, n17690, n17691, n17692, n17693, n17694, n17695, n17696,
         n17697, n17698, n17699, n17700, n17701, n17702, n17703, n17704,
         n17705, n17706, n17707, n17708, n17709, n17710, n17711, n17712,
         n17713, n17714, n17715, n17716, n17717, n17718, n17719, n17720,
         n17721, n17722, n17723, n17724, n17725, n17726, n17727, n17728,
         n17729, n17730, n17731, n17732, n17733, n17734, n17735, n17736,
         n17737, n17738, n17739, n17740, n17741, n17742, n17743, n17744,
         n17745, n17746, n17747, n17748, n17749, n17750, n17751, n17752,
         n17753, n17754, n17755, n17756, n17757, n17758, n17759, n17760,
         n17761, n17762, n17763, n17764, n17765, n17766, n17767, n17768,
         n17769, n17770, n17771, n17772, n17773, n17774, n17775, n17776,
         n17777, n17778, n17779, n17780, n17781, n17782, n17783, n17784,
         n17785, n17786, n17787, n17788, n17789, n17790, n17791, n17792,
         n17793, n17794, n17795, n17796, n17797, n17798, n17799, n17800,
         n17801, n17802, n17803, n17804, n17805, n17806, n17807, n17808,
         n17809, n17810, n17811, n17812, n17813, n17814, n17815, n17816,
         n17817, n17818, n17819, n17820, n17821, n17822, n17823, n17824,
         n17825, n17826, n17827, n17828, n17829, n17830, n17831, n17832,
         n17833, n17834, n17835, n17836, n17837, n17838, n17839, n17840,
         n17841, n17842, n17843, n17844, n17845, n17846, n17847, n17848,
         n17849, n17850, n17851, n17852, n17853, n17854, n17855, n17856,
         n17857, n17858, n17859, n17860, n17861, n17862, n17863, n17864,
         n17865, n17866, n17867, n17868, n17869, n17870, n17871, n17872,
         n17873, n17874, n17875, n17876, n17877, n17878, n17879, n17880,
         n17881, n17882, n17883, n17884, n17885, n17886, n17887, n17888,
         n17889, n17890, n17891, n17892, n17893, n17894, n17895, n17896,
         n17897, n17898, n17899, n17900, n17901, n17902, n17903, n17904,
         n17905, n17906, n17907, n17908, n17909, n17910, n17911, n17912,
         n17913, n17914, n17915, n17916, n17917, n17918, n17919, n17920,
         n17921, n17922, n17923, n17924, n17925, n17926, n17927, n17928,
         n17929, n17930, n17931, n17932, n17933, n17934, n17935, n17936,
         n17937, n17938, n17939, n17940, n17941, n17942, n17943, n17944,
         n17945, n17946, n17947, n17948, n17949, n17950, n17951, n17952,
         n17953, n17954, n17955, n17956, n17957, n17958, n17959, n17960,
         n17961, n17962, n17963, n17964, n17965, n17966, n17967, n17968,
         n17969, n17970, n17971, n17972, n17973, n17974, n17975, n17976,
         n17977, n17978, n17979, n17980, n17981, n17982, n17983, n17984,
         n17985, n17986, n17987, n17988, n17989, n17990, n17991, n17992,
         n17993, n17994, n17995, n17996, n17997, n17998, n17999, n18000,
         n18001, n18002, n18003, n18004, n18005, n18006, n18007, n18008,
         n18009, n18010, n18011, n18012, n18013, n18014, n18015, n18016,
         n18017, n18018, n18019, n18020, n18021, n18022, n18023, n18024,
         n18025, n18026, n18027, n18028, n18029, n18030, n18031, n18032,
         n18033, n18034, n18035, n18036, n18037, n18038, n18039, n18040,
         n18041, n18042, n18043, n18044, n18045, n18046, n18047, n18048,
         n18049, n18050, n18051, n18052, n18053, n18054, n18055, n18056,
         n18057, n18058, n18059, n18060, n18061, n18062, n18063, n18064,
         n18065, n18066, n18067, n18068, n18069, n18070, n18071, n18072,
         n18073, n18074, n18075, n18076, n18077, n18078, n18079, n18080,
         n18081, n18082, n18083, n18084, n18085, n18086, n18087, n18088,
         n18089, n18090, n18091, n18092, n18093, n18094, n18095, n18096,
         n18097, n18098, n18099, n18100, n18101, n18102, n18103, n18104,
         n18105, n18106, n18107, n18108, n18109, n18110, n18111, n18112,
         n18113, n18114, n18115, n18116, n18117, n18118, n18119, n18120,
         n18121, n18122, n18123, n18124, n18125, n18126, n18127, n18128,
         n18129, n18130, n18131, n18132, n18133, n18134, n18135, n18136,
         n18137, n18138, n18139, n18140, n18141, n18142, n18143, n18144,
         n18145, n18146, n18147, n18148, n18149, n18150, n18151, n18152,
         n18153, n18154, n18155, n18156, n18157, n18158, n18159, n18160,
         n18161, n18162, n18163, n18164, n18165, n18166, n18167, n18168,
         n18169, n18170, n18171, n18172, n18173, n18174, n18175, n18176,
         n18177, n18178, n18179, n18180, n18181, n18182, n18183, n18184,
         n18185, n18186, n18187, n18188, n18189, n18190, n18191, n18192,
         n18193, n18194, n18195, n18196, n18197, n18198, n18199, n18200,
         n18201, n18202, n18203, n18204, n18205, n18206, n18207, n18208,
         n18209, n18210, n18211, n18212, n18213, n18214, n18215, n18216,
         n18217, n18218, n18219, n18220, n18221, n18222, n18223, n18224,
         n18225, n18226, n18227, n18228, n18229, n18230, n18231, n18232,
         n18233, n18234, n18235, n18236, n18237, n18238, n18239, n18240,
         n18241, n18242, n18243, n18244, n18245, n18246, n18247, n18248,
         n18249, n18250, n18251, n18252, n18253, n18254, n18255, n18256,
         n18257, n18258, n18259, n18260, n18261, n18262, n18263, n18264,
         n18265, n18266, n18267, n18268, n18269, n18270, n18271, n18272,
         n18273, n18274, n18275, n18276, n18277, n18278, n18279, n18280,
         n18281, n18282, n18283, n18284, n18285, n18286, n18287, n18288,
         n18289, n18290, n18291, n18292, n18293, n18294, n18295, n18296,
         n18297, n18298, n18299, n18300, n18301, n18302, n18303, n18304,
         n18305, n18306, n18307, n18308, n18309, n18310, n18311, n18312,
         n18313, n18314, n18315, n18316, n18317, n18318, n18319, n18320,
         n18321, n18322, n18323, n18324, n18325, n18326, n18327, n18328,
         n18329, n18330, n18331, n18332, n18333, n18334, n18335, n18336,
         n18337, n18338, n18339, n18340, n18341, n18342, n18343, n18344,
         n18345, n18346, n18347, n18348, n18349, n18350, n18351, n18352,
         n18353, n18354, n18355, n18356, n18357, n18358, n18359, n18360,
         n18361, n18362, n18363, n18364, n18365, n18366, n18367, n18368,
         n18369, n18370, n18371, n18372, n18373, n18374, n18375, n18376,
         n18377, n18378, n18379, n18380, n18381, n18382, n18383, n18384,
         n18385, n18386, n18387, n18388, n18389, n18390, n18391, n18392,
         n18393, n18394, n18395, n18396, n18397, n18398, n18399, n18400,
         n18401, n18402, n18403, n18404, n18405, n18406, n18407, n18408,
         n18409, n18410, n18411, n18412, n18413, n18414, n18415, n18416,
         n18417, n18418, n18419, n18420, n18421, n18422, n18423, n18424,
         n18425, n18426, n18427, n18428, n18429, n18430, n18431, n18432,
         n18433, n18434, n18435, n18436, n18437, n18438, n18439, n18440,
         n18441, n18442, n18443, n18444, n18445, n18446, n18447, n18448,
         n18449, n18450, n18451, n18452, n18453, n18454, n18455, n18456,
         n18457, n18458, n18459, n18460, n18461, n18462, n18463, n18464,
         n18465, n18466, n18467, n18468, n18469, n18470, n18471, n18472,
         n18473, n18474, n18475, n18476, n18477, n18478, n18479, n18480,
         n18481, n18482, n18483, n18484, n18485, n18486, n18487, n18488,
         n18489, n18490, n18491, n18492, n18493, n18494, n18495, n18496,
         n18497, n18498, n18499, n18500, n18501, n18502, n18503, n18504,
         n18505, n18506, n18507, n18508, n18509, n18510, n18511, n18512,
         n18513, n18514, n18515, n18516, n18517, n18518, n18519, n18520,
         n18521, n18522, n18523, n18524, n18525, n18526, n18527, n18528,
         n18529, n18530, n18531, n18532, n18533, n18534, n18535, n18536,
         n18537, n18538, n18539, n18540, n18541, n18542, n18543, n18544,
         n18545, n18546, n18547, n18548, n18549, n18550, n18551, n18552,
         n18553, n18554, n18555, n18556, n18557, n18558, n18559, n18560,
         n18561, n18562, n18563, n18564, n18565, n18566, n18567, n18568,
         n18569, n18570, n18571, n18572, n18573, n18574, n18575, n18576,
         n18577, n18578, n18579, n18580, n18581, n18582, n18583, n18584,
         n18585, n18586, n18587, n18588, n18589, n18590, n18591, n18592,
         n18593, n18594, n18595, n18596, n18597, n18598, n18599, n18600,
         n18601, n18602, n18603, n18604, n18605, n18606, n18607, n18608,
         n18609, n18610, n18611, n18612, n18613, n18614, n18615, n18616,
         n18617, n18618, n18619, n18620, n18621, n18622, n18623, n18624,
         n18625, n18626, n18627, n18628, n18629, n18630, n18631, n18632,
         n18633, n18634, n18635, n18636, n18637, n18638, n18639, n18640,
         n18641, n18642, n18643, n18644, n18645, n18646, n18647, n18648,
         n18649, n18650, n18651, n18652, n18653, n18654, n18655, n18656,
         n18657, n18658, n18659, n18660, n18661, n18662, n18663, n18664,
         n18665, n18666, n18667, n18668, n18669, n18670, n18671, n18672,
         n18673, n18674, n18675, n18676, n18677, n18678, n18679, n18680,
         n18681, n18682, n18683, n18684, n18685, n18686, n18687, n18688,
         n18689, n18690, n18691, n18692, n18693, n18694, n18695, n18696,
         n18697, n18698, n18699, n18700, n18701, n18702, n18703, n18704,
         n18705, n18706, n18707, n18708, n18709, n18710, n18711, n18712,
         n18713, n18714, n18715, n18716, n18717, n18718, n18719, n18720,
         n18721, n18722, n18723, n18724, n18725, n18726, n18727, n18728,
         n18729, n18730, n18731, n18732, n18733, n18734, n18735, n18736,
         n18737, n18738, n18739, n18740, n18741, n18742, n18743, n18744,
         n18745, n18746, n18747, n18748, n18749, n18750, n18751, n18752,
         n18753, n18754, n18755, n18756, n18757, n18758, n18759, n18760,
         n18761, n18762, n18763, n18764, n18765, n18766, n18767, n18768,
         n18769, n18770, n18771, n18772, n18773, n18774, n18775, n18776,
         n18777, n18778, n18779, n18780, n18781, n18782, n18783, n18784,
         n18785, n18786, n18787, n18788, n18789, n18790, n18791, n18792,
         n18793, n18794, n18795, n18796, n18797, n18798, n18799, n18800,
         n18801, n18802, n18803, n18804, n18805, n18806, n18807, n18808,
         n18809, n18810, n18811, n18812, n18813, n18814, n18815, n18816,
         n18817, n18818, n18819, n18820, n18821, n18822, n18823, n18824,
         n18825, n18826, n18827, n18828, n18829, n18830, n18831, n18832,
         n18833, n18834, n18835, n18836, n18837, n18838, n18839, n18840,
         n18841, n18842, n18843, n18844, n18845, n18846, n18847, n18848,
         n18849, n18850, n18851, n18852, n18853, n18854, n18855, n18856,
         n18857, n18858, n18859, n18860, n18861, n18862, n18863, n18864,
         n18865, n18866, n18867, n18868, n18869, n18870, n18871, n18872,
         n18873, n18874, n18875, n18876, n18877, n18878, n18879, n18880,
         n18881, n18882, n18883, n18884, n18885, n18886, n18887, n18888,
         n18889, n18890, n18891, n18892, n18893, n18894, n18895, n18896,
         n18897, n18898, n18899, n18900, n18901, n18902, n18903, n18904,
         n18905, n18906, n18907, n18908, n18909, n18910, n18911, n18912,
         n18913, n18914, n18915, n18916, n18917, n18918, n18919, n18920,
         n18921, n18922, n18923, n18924, n18925, n18926, n18927, n18928,
         n18929, n18930, n18931, n18932, n18933, n18934, n18935, n18936,
         n18937, n18938, n18939, n18940, n18941, n18942, n18943, n18944,
         n18945, n18946, n18947, n18948, n18949, n18950, n18951, n18952,
         n18953, n18954, n18955, n18956, n18957, n18958, n18959, n18960,
         n18961, n18962, n18963, n18964, n18965, n18966, n18967, n18968,
         n18969, n18970, n18971, n18972, n18973, n18974, n18975, n18976,
         n18977, n18978, n18979, n18980, n18981, n18982, n18983, n18984,
         n18985, n18986, n18987, n18988, n18989, n18990, n18991, n18992,
         n18993, n18994, n18995, n18996, n18997, n18998, n18999, n19000,
         n19001, n19002, n19003, n19004, n19005, n19006, n19007, n19008,
         n19009, n19010, n19011, n19012, n19013, n19014, n19015, n19016,
         n19017, n19018, n19019, n19020, n19021, n19022, n19023, n19024,
         n19025, n19026, n19027, n19028, n19029, n19030, n19031, n19032,
         n19033, n19034, n19035, n19036, n19037, n19038, n19039, n19040,
         n19041, n19042, n19043, n19044, n19045, n19046, n19047, n19048,
         n19049, n19050, n19051, n19052, n19053, n19054, n19055, n19056,
         n19057, n19058, n19059, n19060, n19061, n19062, n19063, n19064,
         n19065, n19066, n19067, n19068, n19069, n19070, n19071, n19072,
         n19073, n19074, n19075, n19076, n19077, n19078, n19079, n19080,
         n19081, n19082, n19083, n19084, n19085, n19086, n19087, n19088,
         n19089, n19090, n19091, n19092, n19093, n19094, n19095, n19096,
         n19097, n19098, n19099, n19100, n19101, n19102, n19103, n19104,
         n19105, n19106, n19107, n19108, n19109, n19110, n19111, n19112,
         n19113, n19114, n19115, n19116, n19117, n19118, n19119, n19120,
         n19121, n19122, n19123, n19124, n19125, n19126, n19127, n19128,
         n19129, n19130, n19131, n19132, n19133, n19134, n19135, n19136,
         n19137, n19138, n19139, n19140, n19141, n19142, n19143, n19144,
         n19145, n19146, n19147, n19148, n19149, n19150, n19151, n19152,
         n19153, n19154, n19155, n19156, n19157, n19158, n19159, n19160,
         n19161, n19162, n19163, n19164, n19165, n19166, n19167, n19168,
         n19169, n19170, n19171, n19172, n19173, n19174, n19175, n19176,
         n19177, n19178, n19179, n19180, n19181, n19182, n19183, n19184,
         n19185, n19186, n19187, n19188, n19189, n19190, n19191, n19192,
         n19193, n19194, n19195, n19196, n19197, n19198, n19199, n19200,
         n19201, n19202, n19203, n19204, n19205, n19206, n19207, n19208,
         n19209, n19210, n19211, n19212, n19213, n19214, n19215, n19216,
         n19217, n19218, n19219, n19220, n19221, n19222, n19223, n19224,
         n19225, n19226, n19227, n19228, n19229, n19230, n19231, n19232,
         n19233, n19234, n19235, n19236, n19237, n19238, n19239, n19240,
         n19241, n19242, n19243, n19244, n19245, n19246, n19247, n19248,
         n19249, n19250, n19251, n19252, n19253, n19254, n19255, n19256,
         n19257, n19258, n19259, n19260, n19261, n19262, n19263, n19264,
         n19265, n19266, n19267, n19268, n19269, n19270, n19271, n19272,
         n19273, n19274, n19275, n19276, n19277, n19278, n19279, n19280,
         n19281, n19282, n19283, n19284, n19285, n19286, n19287, n19288,
         n19289, n19290, n19291, n19292, n19293, n19294, n19295, n19296,
         n19297, n19298, n19299, n19300, n19301, n19302, n19303, n19304,
         n19305, n19306, n19307, n19308, n19309, n19310, n19311, n19312,
         n19313, n19314, n19315, n19316, n19317, n19318, n19319, n19320,
         n19321, n19322, n19323, n19324, n19325, n19326, n19327, n19328,
         n19329, n19330, n19331, n19332, n19333, n19334, n19335, n19336,
         n19337, n19338, n19339, n19340, n19341, n19342, n19343, n19344,
         n19345, n19346, n19347, n19348, n19349, n19350, n19351, n19352,
         n19353, n19354, n19355, n19356, n19357, n19358, n19359, n19360,
         n19361, n19362, n19363, n19364, n19365, n19366, n19367, n19368,
         n19369, n19370, n19371, n19372, n19373, n19374, n19375, n19376,
         n19377, n19378, n19379, n19380, n19381, n19382, n19383, n19384,
         n19385, n19386, n19387, n19388, n19389, n19390, n19391, n19392,
         n19393, n19394, n19395, n19396, n19397, n19398, n19399, n19400,
         n19401, n19402, n19403, n19404, n19405, n19406, n19407, n19408,
         n19409, n19410, n19411, n19412, n19413, n19414, n19415, n19416,
         n19417, n19418, n19419, n19420, n19421, n19422, n19423, n19424,
         n19425, n19426, n19427, n19428, n19429, n19430, n19431, n19432,
         n19433, n19434, n19435, n19436, n19437, n19438, n19439, n19440,
         n19441, n19442, n19443, n19444, n19445, n19446, n19447, n19448,
         n19449, n19450, n19451, n19452, n19453, n19454, n19455, n19456,
         n19457, n19458, n19459, n19460, n19461, n19462, n19463, n19464,
         n19465, n19466, n19467, n19468, n19469, n19470, n19471, n19472,
         n19473, n19474, n19475, n19476, n19477, n19478, n19479, n19480,
         n19481, n19482, n19483, n19484, n19485, n19486, n19487, n19488,
         n19489, n19490, n19491, n19492, n19493, n19494, n19495, n19496,
         n19497, n19498, n19499, n19500, n19501, n19502, n19503, n19504,
         n19505, n19506, n19507, n19508, n19509, n19510, n19511, n19512,
         n19513, n19514, n19515, n19516, n19517, n19518, n19519, n19520,
         n19521, n19522, n19523, n19524, n19525, n19526, n19527, n19528,
         n19529, n19530, n19531, n19532, n19533, n19534, n19535, n19536,
         n19537, n19538, n19539, n19540, n19541, n19542, n19543, n19544,
         n19545, n19546, n19547, n19548, n19549, n19550, n19551, n19552,
         n19553, n19554, n19555, n19556, n19557, n19558, n19559, n19560,
         n19561, n19562, n19563, n19564, n19565, n19566, n19567, n19568,
         n19569, n19570, n19571, n19572, n19573, n19574, n19575, n19576,
         n19577, n19578, n19579, n19580, n19581, n19582, n19583, n19584,
         n19585, n19586, n19587, n19588, n19589, n19590, n19591, n19592,
         n19593, n19594, n19595, n19596, n19597, n19598, n19599, n19600,
         n19601, n19602, n19603, n19604, n19605, n19606, n19607, n19608,
         n19609, n19610, n19611, n19612, n19613, n19614, n19615, n19616,
         n19617, n19618, n19619, n19620, n19621, n19622, n19623, n19624,
         n19625, n19626, n19627, n19628, n19629, n19630, n19631, n19632,
         n19633, n19634, n19635, n19636, n19637, n19638, n19639, n19640,
         n19641, n19642, n19643, n19644, n19645, n19646, n19647, n19648,
         n19649, n19650, n19651, n19652, n19653, n19654, n19655, n19656,
         n19657, n19658, n19659, n19660, n19661, n19662, n19663, n19664,
         n19665, n19666, n19667, n19668, n19669, n19670, n19671, n19672,
         n19673, n19674, n19675, n19676, n19677, n19678, n19679, n19680,
         n19681, n19682, n19683, n19684, n19685, n19686, n19687, n19688,
         n19689, n19690, n19691, n19692, n19693, n19694, n19695, n19696,
         n19697, n19698, n19699, n19700, n19701, n19702, n19703, n19704,
         n19705, n19706, n19707, n19708, n19709, n19710, n19711, n19712,
         n19713, n19714, n19715, n19716, n19717, n19718, n19719, n19720,
         n19721, n19722, n19723, n19724, n19725, n19726, n19727, n19728,
         n19729, n19730, n19731, n19732, n19733, n19734, n19735, n19736,
         n19737, n19738, n19739, n19740, n19741, n19742, n19743, n19744,
         n19745, n19746, n19747, n19748, n19749, n19750, n19751, n19752,
         n19753, n19754, n19755, n19756, n19757, n19758, n19759, n19760,
         n19761, n19762, n19763, n19764, n19765, n19766, n19767, n19768,
         n19769, n19770, n19771, n19772, n19773, n19774, n19775, n19776,
         n19777, n19778, n19779, n19780, n19781, n19782, n19783, n19784,
         n19785, n19786, n19787, n19788, n19789, n19790, n19791, n19792,
         n19793, n19794, n19795, n19796, n19797, n19798, n19799, n19800,
         n19801, n19802, n19803, n19804, n19805, n19806, n19807, n19808,
         n19809, n19810, n19811, n19812, n19813, n19814, n19815, n19816,
         n19817, n19818, n19819, n19820, n19821, n19822, n19823, n19824,
         n19825, n19826, n19827, n19828, n19829, n19830, n19831, n19832,
         n19833, n19834, n19835, n19836, n19837, n19838, n19839, n19840,
         n19841, n19842, n19843, n19844, n19845, n19846, n19847, n19848,
         n19849, n19850, n19851, n19852, n19853, n19854, n19855, n19856,
         n19857, n19858, n19859, n19860, n19861, n19862, n19863, n19864,
         n19865, n19866, n19867, n19868, n19869, n19870, n19871, n19872,
         n19873, n19874, n19875, n19876, n19877, n19878, n19879, n19880,
         n19881, n19882, n19883, n19884, n19885, n19886, n19887, n19888,
         n19889, n19890, n19891, n19892, n19893, n19894, n19895, n19896,
         n19897, n19898, n19899, n19900, n19901, n19902, n19903, n19904,
         n19905, n19906, n19907, n19908, n19909, n19910, n19911, n19912;
  assign \MULT3/B__[0]  = e_input[0];

  IV U2 ( .A(n16747), .Z(n19720) );
  ANDN U3 ( .A(n2), .B(n3), .Z(o) );
  NANDN U4 ( .B(n3), .A(n4), .Z(n2) );
  XOR U5 ( .A(n5), .B(n6), .Z(n4) );
  AND U6 ( .A(n7), .B(n8), .Z(n5) );
  XOR U7 ( .A(n9), .B(n10), .Z(n8) );
  XNOR U8 ( .A(n11), .B(n6), .Z(n7) );
  XOR U9 ( .A(n12), .B(n13), .Z(n6) );
  ANDN U10 ( .A(n14), .B(n15), .Z(n13) );
  XNOR U11 ( .A(n9), .B(n12), .Z(n14) );
  NANDN U12 ( .B(n16), .A(n17), .Z(n3) );
  OR U13 ( .A(n11), .B(n16), .Z(n17) );
  XOR U14 ( .A(n18), .B(n9), .Z(n11) );
  IV U15 ( .A(n15), .Z(n18) );
  XOR U16 ( .A(n12), .B(n10), .Z(n15) );
  XNOR U17 ( .A(n19), .B(n20), .Z(n10) );
  AND U18 ( .A(n21), .B(n22), .Z(n20) );
  XNOR U19 ( .A(n19), .B(n23), .Z(n22) );
  XOR U20 ( .A(n24), .B(n25), .Z(n12) );
  AND U21 ( .A(n26), .B(n27), .Z(n25) );
  XNOR U22 ( .A(n9), .B(n24), .Z(n27) );
  NANDN U23 ( .B(n28), .A(n29), .Z(n16) );
  NANDN U24 ( .B(n28), .A(n30), .Z(n29) );
  XNOR U25 ( .A(n9), .B(n26), .Z(n30) );
  XOR U26 ( .A(n31), .B(n23), .Z(n26) );
  XNOR U27 ( .A(n32), .B(n33), .Z(n23) );
  ANDN U28 ( .A(n34), .B(n35), .Z(n33) );
  XNOR U29 ( .A(n32), .B(n36), .Z(n34) );
  XNOR U30 ( .A(n21), .B(n24), .Z(n31) );
  XOR U31 ( .A(n37), .B(n38), .Z(n24) );
  AND U32 ( .A(n39), .B(n40), .Z(n38) );
  XNOR U33 ( .A(n9), .B(n37), .Z(n40) );
  XOR U34 ( .A(n19), .B(n41), .Z(n21) );
  ANDN U35 ( .A(n42), .B(n43), .Z(n41) );
  XOR U36 ( .A(n44), .B(n45), .Z(n19) );
  AND U37 ( .A(n46), .B(n47), .Z(n45) );
  XNOR U38 ( .A(n44), .B(n48), .Z(n47) );
  NANDN U39 ( .B(n49), .A(n50), .Z(n28) );
  NANDN U40 ( .B(n49), .A(n51), .Z(n50) );
  XNOR U41 ( .A(n9), .B(n39), .Z(n51) );
  XOR U42 ( .A(n52), .B(n48), .Z(n39) );
  XOR U43 ( .A(n36), .B(n53), .Z(n48) );
  IV U44 ( .A(n35), .Z(n53) );
  XNOR U45 ( .A(n32), .B(n54), .Z(n35) );
  AND U46 ( .A(n42), .B(n80), .Z(n54) );
  XOR U47 ( .A(n55), .B(n56), .Z(n32) );
  ANDN U48 ( .A(n57), .B(n58), .Z(n56) );
  XNOR U49 ( .A(n55), .B(n59), .Z(n57) );
  XNOR U50 ( .A(n60), .B(n61), .Z(n36) );
  ANDN U51 ( .A(n62), .B(n63), .Z(n61) );
  XNOR U52 ( .A(n60), .B(n64), .Z(n62) );
  XNOR U53 ( .A(n46), .B(n37), .Z(n52) );
  XOR U54 ( .A(n65), .B(n66), .Z(n37) );
  AND U55 ( .A(n67), .B(n68), .Z(n66) );
  XNOR U56 ( .A(n9), .B(n65), .Z(n68) );
  XOR U57 ( .A(n44), .B(n69), .Z(n46) );
  ANDN U58 ( .A(n80), .B(n43), .Z(n69) );
  XOR U59 ( .A(n70), .B(n71), .Z(n44) );
  AND U60 ( .A(n72), .B(n73), .Z(n71) );
  XNOR U61 ( .A(n70), .B(n74), .Z(n73) );
  NANDN U62 ( .B(n75), .A(n76), .Z(n49) );
  NANDN U63 ( .B(n75), .A(n77), .Z(n76) );
  XNOR U64 ( .A(n9), .B(n67), .Z(n77) );
  XOR U65 ( .A(n78), .B(n74), .Z(n67) );
  XOR U66 ( .A(n59), .B(n79), .Z(n74) );
  IV U67 ( .A(n58), .Z(n79) );
  XNOR U68 ( .A(n55), .B(n80), .Z(n58) );
  XOR U69 ( .A(n81), .B(n82), .Z(n55) );
  ANDN U70 ( .A(n83), .B(n84), .Z(n82) );
  XNOR U71 ( .A(n81), .B(n85), .Z(n83) );
  XOR U72 ( .A(n64), .B(n86), .Z(n59) );
  IV U73 ( .A(n63), .Z(n86) );
  XNOR U74 ( .A(n60), .B(n87), .Z(n63) );
  AND U75 ( .A(n42), .B(n159), .Z(n87) );
  XOR U76 ( .A(n88), .B(n89), .Z(n60) );
  ANDN U77 ( .A(n90), .B(n91), .Z(n89) );
  XNOR U78 ( .A(n88), .B(n92), .Z(n90) );
  XNOR U79 ( .A(n93), .B(n94), .Z(n64) );
  ANDN U80 ( .A(n95), .B(n96), .Z(n94) );
  XNOR U81 ( .A(n93), .B(n97), .Z(n95) );
  XNOR U82 ( .A(n72), .B(n65), .Z(n78) );
  XOR U83 ( .A(n98), .B(n99), .Z(n65) );
  AND U84 ( .A(n100), .B(n101), .Z(n99) );
  XNOR U85 ( .A(n9), .B(n98), .Z(n101) );
  XOR U86 ( .A(n70), .B(n102), .Z(n72) );
  ANDN U87 ( .A(n159), .B(n43), .Z(n102) );
  XOR U88 ( .A(n103), .B(n104), .Z(n70) );
  AND U89 ( .A(n105), .B(n106), .Z(n104) );
  XNOR U90 ( .A(n103), .B(n107), .Z(n106) );
  NANDN U91 ( .B(n108), .A(n109), .Z(n75) );
  NANDN U92 ( .B(n108), .A(n110), .Z(n109) );
  XNOR U93 ( .A(n9), .B(n100), .Z(n110) );
  XOR U94 ( .A(n111), .B(n107), .Z(n100) );
  XOR U95 ( .A(n85), .B(n112), .Z(n107) );
  IV U96 ( .A(n84), .Z(n112) );
  XNOR U97 ( .A(n81), .B(n113), .Z(n84) );
  XOR U98 ( .A(n114), .B(n115), .Z(n81) );
  ANDN U99 ( .A(n116), .B(n117), .Z(n115) );
  XNOR U100 ( .A(n114), .B(n118), .Z(n116) );
  XOR U101 ( .A(n92), .B(n119), .Z(n85) );
  IV U102 ( .A(n91), .Z(n119) );
  XNOR U103 ( .A(n88), .B(n113), .Z(n91) );
  AND U104 ( .A(n159), .B(n80), .Z(n113) );
  XOR U105 ( .A(n120), .B(n121), .Z(n88) );
  ANDN U106 ( .A(n122), .B(n123), .Z(n121) );
  XNOR U107 ( .A(n120), .B(n124), .Z(n122) );
  XOR U108 ( .A(n97), .B(n125), .Z(n92) );
  IV U109 ( .A(n96), .Z(n125) );
  XNOR U110 ( .A(n93), .B(n126), .Z(n96) );
  AND U111 ( .A(n42), .B(n264), .Z(n126) );
  XOR U112 ( .A(n127), .B(n128), .Z(n93) );
  ANDN U113 ( .A(n129), .B(n130), .Z(n128) );
  XNOR U114 ( .A(n127), .B(n131), .Z(n129) );
  XNOR U115 ( .A(n132), .B(n133), .Z(n97) );
  ANDN U116 ( .A(n134), .B(n135), .Z(n133) );
  XNOR U117 ( .A(n132), .B(n136), .Z(n134) );
  XNOR U118 ( .A(n105), .B(n98), .Z(n111) );
  XOR U119 ( .A(n137), .B(n138), .Z(n98) );
  AND U120 ( .A(n139), .B(n140), .Z(n138) );
  XNOR U121 ( .A(n9), .B(n137), .Z(n140) );
  XOR U122 ( .A(n103), .B(n141), .Z(n105) );
  ANDN U123 ( .A(n264), .B(n43), .Z(n141) );
  XOR U124 ( .A(n142), .B(n143), .Z(n103) );
  AND U125 ( .A(n144), .B(n145), .Z(n143) );
  XNOR U126 ( .A(n142), .B(n146), .Z(n145) );
  NANDN U127 ( .B(n147), .A(n148), .Z(n108) );
  NANDN U128 ( .B(n147), .A(n149), .Z(n148) );
  XNOR U129 ( .A(n9), .B(n139), .Z(n149) );
  XOR U130 ( .A(n150), .B(n146), .Z(n139) );
  XOR U131 ( .A(n118), .B(n151), .Z(n146) );
  IV U132 ( .A(n117), .Z(n151) );
  XNOR U133 ( .A(n114), .B(n152), .Z(n117) );
  XOR U134 ( .A(n153), .B(n154), .Z(n114) );
  ANDN U135 ( .A(n155), .B(n156), .Z(n154) );
  XNOR U136 ( .A(n153), .B(n157), .Z(n155) );
  XOR U137 ( .A(n124), .B(n158), .Z(n118) );
  IV U138 ( .A(n123), .Z(n158) );
  XNOR U139 ( .A(n120), .B(n159), .Z(n123) );
  XOR U140 ( .A(n160), .B(n161), .Z(n120) );
  ANDN U141 ( .A(n162), .B(n163), .Z(n161) );
  XNOR U142 ( .A(n160), .B(n164), .Z(n162) );
  XOR U143 ( .A(n131), .B(n165), .Z(n124) );
  IV U144 ( .A(n130), .Z(n165) );
  XNOR U145 ( .A(n127), .B(n152), .Z(n130) );
  AND U146 ( .A(n264), .B(n80), .Z(n152) );
  XOR U147 ( .A(n166), .B(n167), .Z(n127) );
  ANDN U148 ( .A(n168), .B(n169), .Z(n167) );
  XNOR U149 ( .A(n166), .B(n170), .Z(n168) );
  XOR U150 ( .A(n136), .B(n171), .Z(n131) );
  IV U151 ( .A(n135), .Z(n171) );
  XNOR U152 ( .A(n132), .B(n172), .Z(n135) );
  AND U153 ( .A(n42), .B(n395), .Z(n172) );
  XOR U154 ( .A(n173), .B(n174), .Z(n132) );
  ANDN U155 ( .A(n175), .B(n176), .Z(n174) );
  XNOR U156 ( .A(n173), .B(n177), .Z(n175) );
  XNOR U157 ( .A(n178), .B(n179), .Z(n136) );
  ANDN U158 ( .A(n180), .B(n181), .Z(n179) );
  XNOR U159 ( .A(n178), .B(n182), .Z(n180) );
  XNOR U160 ( .A(n144), .B(n137), .Z(n150) );
  XOR U161 ( .A(n183), .B(n184), .Z(n137) );
  AND U162 ( .A(n185), .B(n186), .Z(n184) );
  XNOR U163 ( .A(n9), .B(n183), .Z(n186) );
  XOR U164 ( .A(n142), .B(n187), .Z(n144) );
  ANDN U165 ( .A(n395), .B(n43), .Z(n187) );
  XOR U166 ( .A(n188), .B(n189), .Z(n142) );
  AND U167 ( .A(n190), .B(n191), .Z(n189) );
  XNOR U168 ( .A(n188), .B(n192), .Z(n191) );
  NANDN U169 ( .B(n193), .A(n194), .Z(n147) );
  NANDN U170 ( .B(n193), .A(n195), .Z(n194) );
  XNOR U171 ( .A(n9), .B(n185), .Z(n195) );
  XOR U172 ( .A(n196), .B(n192), .Z(n185) );
  XOR U173 ( .A(n157), .B(n197), .Z(n192) );
  IV U174 ( .A(n156), .Z(n197) );
  XNOR U175 ( .A(n153), .B(n198), .Z(n156) );
  XOR U176 ( .A(n199), .B(n200), .Z(n153) );
  ANDN U177 ( .A(n201), .B(n202), .Z(n200) );
  XNOR U178 ( .A(n199), .B(n203), .Z(n201) );
  XOR U179 ( .A(n164), .B(n204), .Z(n157) );
  IV U180 ( .A(n163), .Z(n204) );
  XNOR U181 ( .A(n160), .B(n205), .Z(n163) );
  XOR U182 ( .A(n206), .B(n207), .Z(n160) );
  ANDN U183 ( .A(n208), .B(n209), .Z(n207) );
  XNOR U184 ( .A(n206), .B(n210), .Z(n208) );
  XOR U185 ( .A(n170), .B(n211), .Z(n164) );
  IV U186 ( .A(n169), .Z(n211) );
  XNOR U187 ( .A(n166), .B(n205), .Z(n169) );
  AND U188 ( .A(n264), .B(n159), .Z(n205) );
  XOR U189 ( .A(n212), .B(n213), .Z(n166) );
  ANDN U190 ( .A(n214), .B(n215), .Z(n213) );
  XNOR U191 ( .A(n212), .B(n216), .Z(n214) );
  XOR U192 ( .A(n177), .B(n217), .Z(n170) );
  IV U193 ( .A(n176), .Z(n217) );
  XNOR U194 ( .A(n173), .B(n198), .Z(n176) );
  AND U195 ( .A(n395), .B(n80), .Z(n198) );
  XOR U196 ( .A(n218), .B(n219), .Z(n173) );
  ANDN U197 ( .A(n220), .B(n221), .Z(n219) );
  XNOR U198 ( .A(n218), .B(n222), .Z(n220) );
  XOR U199 ( .A(n182), .B(n223), .Z(n177) );
  IV U200 ( .A(n181), .Z(n223) );
  XNOR U201 ( .A(n178), .B(n224), .Z(n181) );
  AND U202 ( .A(n42), .B(n552), .Z(n224) );
  XOR U203 ( .A(n225), .B(n226), .Z(n178) );
  ANDN U204 ( .A(n227), .B(n228), .Z(n226) );
  XNOR U205 ( .A(n225), .B(n229), .Z(n227) );
  XNOR U206 ( .A(n230), .B(n231), .Z(n182) );
  ANDN U207 ( .A(n232), .B(n233), .Z(n231) );
  XNOR U208 ( .A(n230), .B(n234), .Z(n232) );
  XNOR U209 ( .A(n190), .B(n183), .Z(n196) );
  XOR U210 ( .A(n235), .B(n236), .Z(n183) );
  AND U211 ( .A(n237), .B(n238), .Z(n236) );
  XNOR U212 ( .A(n9), .B(n235), .Z(n238) );
  XOR U213 ( .A(n188), .B(n239), .Z(n190) );
  ANDN U214 ( .A(n552), .B(n43), .Z(n239) );
  XOR U215 ( .A(n240), .B(n241), .Z(n188) );
  AND U216 ( .A(n242), .B(n243), .Z(n241) );
  XNOR U217 ( .A(n240), .B(n244), .Z(n243) );
  NANDN U218 ( .B(n245), .A(n246), .Z(n193) );
  NANDN U219 ( .B(n245), .A(n247), .Z(n246) );
  XNOR U220 ( .A(n9), .B(n237), .Z(n247) );
  XOR U221 ( .A(n248), .B(n244), .Z(n237) );
  XOR U222 ( .A(n203), .B(n249), .Z(n244) );
  IV U223 ( .A(n202), .Z(n249) );
  XNOR U224 ( .A(n199), .B(n250), .Z(n202) );
  XOR U225 ( .A(n251), .B(n252), .Z(n199) );
  ANDN U226 ( .A(n253), .B(n254), .Z(n252) );
  XNOR U227 ( .A(n251), .B(n255), .Z(n253) );
  XOR U228 ( .A(n210), .B(n256), .Z(n203) );
  IV U229 ( .A(n209), .Z(n256) );
  XNOR U230 ( .A(n206), .B(n257), .Z(n209) );
  XOR U231 ( .A(n258), .B(n259), .Z(n206) );
  ANDN U232 ( .A(n260), .B(n261), .Z(n259) );
  XNOR U233 ( .A(n258), .B(n262), .Z(n260) );
  XOR U234 ( .A(n216), .B(n263), .Z(n210) );
  IV U235 ( .A(n215), .Z(n263) );
  XNOR U236 ( .A(n212), .B(n264), .Z(n215) );
  XOR U237 ( .A(n265), .B(n266), .Z(n212) );
  ANDN U238 ( .A(n267), .B(n268), .Z(n266) );
  XNOR U239 ( .A(n265), .B(n269), .Z(n267) );
  XOR U240 ( .A(n222), .B(n270), .Z(n216) );
  IV U241 ( .A(n221), .Z(n270) );
  XNOR U242 ( .A(n218), .B(n257), .Z(n221) );
  AND U243 ( .A(n395), .B(n159), .Z(n257) );
  XOR U244 ( .A(n271), .B(n272), .Z(n218) );
  ANDN U245 ( .A(n273), .B(n274), .Z(n272) );
  XNOR U246 ( .A(n271), .B(n275), .Z(n273) );
  XOR U247 ( .A(n229), .B(n276), .Z(n222) );
  IV U248 ( .A(n228), .Z(n276) );
  XNOR U249 ( .A(n225), .B(n250), .Z(n228) );
  AND U250 ( .A(n552), .B(n80), .Z(n250) );
  XOR U251 ( .A(n277), .B(n278), .Z(n225) );
  ANDN U252 ( .A(n279), .B(n280), .Z(n278) );
  XNOR U253 ( .A(n277), .B(n281), .Z(n279) );
  XOR U254 ( .A(n234), .B(n282), .Z(n229) );
  IV U255 ( .A(n233), .Z(n282) );
  XNOR U256 ( .A(n230), .B(n283), .Z(n233) );
  AND U257 ( .A(n42), .B(n736), .Z(n283) );
  XOR U258 ( .A(n284), .B(n285), .Z(n230) );
  ANDN U259 ( .A(n286), .B(n287), .Z(n285) );
  XNOR U260 ( .A(n284), .B(n288), .Z(n286) );
  XNOR U261 ( .A(n289), .B(n290), .Z(n234) );
  ANDN U262 ( .A(n291), .B(n292), .Z(n290) );
  XNOR U263 ( .A(n289), .B(n293), .Z(n291) );
  XNOR U264 ( .A(n242), .B(n235), .Z(n248) );
  XOR U265 ( .A(n294), .B(n295), .Z(n235) );
  AND U266 ( .A(n296), .B(n297), .Z(n295) );
  XNOR U267 ( .A(n9), .B(n294), .Z(n297) );
  XOR U268 ( .A(n240), .B(n298), .Z(n242) );
  ANDN U269 ( .A(n736), .B(n43), .Z(n298) );
  XOR U270 ( .A(n299), .B(n300), .Z(n240) );
  AND U271 ( .A(n301), .B(n302), .Z(n300) );
  XNOR U272 ( .A(n299), .B(n303), .Z(n302) );
  NANDN U273 ( .B(n304), .A(n305), .Z(n245) );
  NANDN U274 ( .B(n304), .A(n306), .Z(n305) );
  XNOR U275 ( .A(n9), .B(n296), .Z(n306) );
  XOR U276 ( .A(n307), .B(n303), .Z(n296) );
  XOR U277 ( .A(n255), .B(n308), .Z(n303) );
  IV U278 ( .A(n254), .Z(n308) );
  XNOR U279 ( .A(n251), .B(n309), .Z(n254) );
  XOR U280 ( .A(n310), .B(n311), .Z(n251) );
  ANDN U281 ( .A(n312), .B(n313), .Z(n311) );
  XNOR U282 ( .A(n310), .B(n314), .Z(n312) );
  XOR U283 ( .A(n262), .B(n315), .Z(n255) );
  IV U284 ( .A(n261), .Z(n315) );
  XNOR U285 ( .A(n258), .B(n316), .Z(n261) );
  XOR U286 ( .A(n317), .B(n318), .Z(n258) );
  ANDN U287 ( .A(n319), .B(n320), .Z(n318) );
  XNOR U288 ( .A(n317), .B(n321), .Z(n319) );
  XOR U289 ( .A(n269), .B(n322), .Z(n262) );
  IV U290 ( .A(n268), .Z(n322) );
  XNOR U291 ( .A(n265), .B(n323), .Z(n268) );
  XOR U292 ( .A(n324), .B(n325), .Z(n265) );
  ANDN U293 ( .A(n326), .B(n327), .Z(n325) );
  XNOR U294 ( .A(n324), .B(n328), .Z(n326) );
  XOR U295 ( .A(n275), .B(n329), .Z(n269) );
  IV U296 ( .A(n274), .Z(n329) );
  XNOR U297 ( .A(n271), .B(n323), .Z(n274) );
  AND U298 ( .A(n395), .B(n264), .Z(n323) );
  XOR U299 ( .A(n330), .B(n331), .Z(n271) );
  ANDN U300 ( .A(n332), .B(n333), .Z(n331) );
  XNOR U301 ( .A(n330), .B(n334), .Z(n332) );
  XOR U302 ( .A(n281), .B(n335), .Z(n275) );
  IV U303 ( .A(n280), .Z(n335) );
  XNOR U304 ( .A(n277), .B(n316), .Z(n280) );
  AND U305 ( .A(n552), .B(n159), .Z(n316) );
  XOR U306 ( .A(n336), .B(n337), .Z(n277) );
  ANDN U307 ( .A(n338), .B(n339), .Z(n337) );
  XNOR U308 ( .A(n336), .B(n340), .Z(n338) );
  XOR U309 ( .A(n288), .B(n341), .Z(n281) );
  IV U310 ( .A(n287), .Z(n341) );
  XNOR U311 ( .A(n284), .B(n309), .Z(n287) );
  AND U312 ( .A(n736), .B(n80), .Z(n309) );
  XOR U313 ( .A(n342), .B(n343), .Z(n284) );
  ANDN U314 ( .A(n344), .B(n345), .Z(n343) );
  XNOR U315 ( .A(n342), .B(n346), .Z(n344) );
  XOR U316 ( .A(n293), .B(n347), .Z(n288) );
  IV U317 ( .A(n292), .Z(n347) );
  XNOR U318 ( .A(n289), .B(n348), .Z(n292) );
  AND U319 ( .A(n42), .B(n948), .Z(n348) );
  XOR U320 ( .A(n349), .B(n350), .Z(n289) );
  ANDN U321 ( .A(n351), .B(n352), .Z(n350) );
  XNOR U322 ( .A(n349), .B(n353), .Z(n351) );
  XNOR U323 ( .A(n354), .B(n355), .Z(n293) );
  ANDN U324 ( .A(n356), .B(n357), .Z(n355) );
  XNOR U325 ( .A(n354), .B(n358), .Z(n356) );
  XNOR U326 ( .A(n301), .B(n294), .Z(n307) );
  XOR U327 ( .A(n359), .B(n360), .Z(n294) );
  AND U328 ( .A(n361), .B(n362), .Z(n360) );
  XNOR U329 ( .A(n9), .B(n359), .Z(n362) );
  XOR U330 ( .A(n299), .B(n363), .Z(n301) );
  ANDN U331 ( .A(n948), .B(n43), .Z(n363) );
  XOR U332 ( .A(n364), .B(n365), .Z(n299) );
  AND U333 ( .A(n366), .B(n367), .Z(n365) );
  XNOR U334 ( .A(n364), .B(n368), .Z(n367) );
  NANDN U335 ( .B(n369), .A(n370), .Z(n304) );
  NANDN U336 ( .B(n369), .A(n371), .Z(n370) );
  XNOR U337 ( .A(n9), .B(n361), .Z(n371) );
  XOR U338 ( .A(n372), .B(n368), .Z(n361) );
  XOR U339 ( .A(n314), .B(n373), .Z(n368) );
  IV U340 ( .A(n313), .Z(n373) );
  XNOR U341 ( .A(n310), .B(n374), .Z(n313) );
  XOR U342 ( .A(n375), .B(n376), .Z(n310) );
  ANDN U343 ( .A(n377), .B(n378), .Z(n376) );
  XNOR U344 ( .A(n375), .B(n379), .Z(n377) );
  XOR U345 ( .A(n321), .B(n380), .Z(n314) );
  IV U346 ( .A(n320), .Z(n380) );
  XNOR U347 ( .A(n317), .B(n381), .Z(n320) );
  XOR U348 ( .A(n382), .B(n383), .Z(n317) );
  ANDN U349 ( .A(n384), .B(n385), .Z(n383) );
  XNOR U350 ( .A(n382), .B(n386), .Z(n384) );
  XOR U351 ( .A(n328), .B(n387), .Z(n321) );
  IV U352 ( .A(n327), .Z(n387) );
  XNOR U353 ( .A(n324), .B(n388), .Z(n327) );
  XOR U354 ( .A(n389), .B(n390), .Z(n324) );
  ANDN U355 ( .A(n391), .B(n392), .Z(n390) );
  XNOR U356 ( .A(n389), .B(n393), .Z(n391) );
  XOR U357 ( .A(n334), .B(n394), .Z(n328) );
  IV U358 ( .A(n333), .Z(n394) );
  XNOR U359 ( .A(n330), .B(n395), .Z(n333) );
  XOR U360 ( .A(n396), .B(n397), .Z(n330) );
  ANDN U361 ( .A(n398), .B(n399), .Z(n397) );
  XNOR U362 ( .A(n396), .B(n400), .Z(n398) );
  XOR U363 ( .A(n340), .B(n401), .Z(n334) );
  IV U364 ( .A(n339), .Z(n401) );
  XNOR U365 ( .A(n336), .B(n388), .Z(n339) );
  AND U366 ( .A(n552), .B(n264), .Z(n388) );
  XOR U367 ( .A(n402), .B(n403), .Z(n336) );
  ANDN U368 ( .A(n404), .B(n405), .Z(n403) );
  XNOR U369 ( .A(n402), .B(n406), .Z(n404) );
  XOR U370 ( .A(n346), .B(n407), .Z(n340) );
  IV U371 ( .A(n345), .Z(n407) );
  XNOR U372 ( .A(n342), .B(n381), .Z(n345) );
  AND U373 ( .A(n736), .B(n159), .Z(n381) );
  XOR U374 ( .A(n408), .B(n409), .Z(n342) );
  ANDN U375 ( .A(n410), .B(n411), .Z(n409) );
  XNOR U376 ( .A(n408), .B(n412), .Z(n410) );
  XOR U377 ( .A(n353), .B(n413), .Z(n346) );
  IV U378 ( .A(n352), .Z(n413) );
  XNOR U379 ( .A(n349), .B(n374), .Z(n352) );
  AND U380 ( .A(n948), .B(n80), .Z(n374) );
  XOR U381 ( .A(n414), .B(n415), .Z(n349) );
  ANDN U382 ( .A(n416), .B(n417), .Z(n415) );
  XNOR U383 ( .A(n414), .B(n418), .Z(n416) );
  XOR U384 ( .A(n358), .B(n419), .Z(n353) );
  IV U385 ( .A(n357), .Z(n419) );
  XNOR U386 ( .A(n354), .B(n420), .Z(n357) );
  AND U387 ( .A(n42), .B(n1185), .Z(n420) );
  XOR U388 ( .A(n421), .B(n422), .Z(n354) );
  ANDN U389 ( .A(n423), .B(n424), .Z(n422) );
  XNOR U390 ( .A(n421), .B(n425), .Z(n423) );
  XNOR U391 ( .A(n426), .B(n427), .Z(n358) );
  ANDN U392 ( .A(n428), .B(n429), .Z(n427) );
  XNOR U393 ( .A(n426), .B(n430), .Z(n428) );
  XNOR U394 ( .A(n366), .B(n359), .Z(n372) );
  XOR U395 ( .A(n431), .B(n432), .Z(n359) );
  AND U396 ( .A(n433), .B(n434), .Z(n432) );
  XNOR U397 ( .A(n9), .B(n431), .Z(n434) );
  XOR U398 ( .A(n364), .B(n435), .Z(n366) );
  ANDN U399 ( .A(n1185), .B(n43), .Z(n435) );
  XOR U400 ( .A(n436), .B(n437), .Z(n364) );
  AND U401 ( .A(n438), .B(n439), .Z(n437) );
  XNOR U402 ( .A(n436), .B(n440), .Z(n439) );
  NANDN U403 ( .B(n441), .A(n442), .Z(n369) );
  NANDN U404 ( .B(n441), .A(n443), .Z(n442) );
  XNOR U405 ( .A(n9), .B(n433), .Z(n443) );
  XOR U406 ( .A(n444), .B(n440), .Z(n433) );
  XOR U407 ( .A(n379), .B(n445), .Z(n440) );
  IV U408 ( .A(n378), .Z(n445) );
  XNOR U409 ( .A(n375), .B(n446), .Z(n378) );
  XOR U410 ( .A(n447), .B(n448), .Z(n375) );
  ANDN U411 ( .A(n449), .B(n450), .Z(n448) );
  XNOR U412 ( .A(n447), .B(n451), .Z(n449) );
  XOR U413 ( .A(n386), .B(n452), .Z(n379) );
  IV U414 ( .A(n385), .Z(n452) );
  XNOR U415 ( .A(n382), .B(n453), .Z(n385) );
  XOR U416 ( .A(n454), .B(n455), .Z(n382) );
  ANDN U417 ( .A(n456), .B(n457), .Z(n455) );
  XNOR U418 ( .A(n454), .B(n458), .Z(n456) );
  XOR U419 ( .A(n393), .B(n459), .Z(n386) );
  IV U420 ( .A(n392), .Z(n459) );
  XNOR U421 ( .A(n389), .B(n460), .Z(n392) );
  XOR U422 ( .A(n461), .B(n462), .Z(n389) );
  ANDN U423 ( .A(n463), .B(n464), .Z(n462) );
  XNOR U424 ( .A(n461), .B(n465), .Z(n463) );
  XOR U425 ( .A(n400), .B(n466), .Z(n393) );
  IV U426 ( .A(n399), .Z(n466) );
  XNOR U427 ( .A(n396), .B(n467), .Z(n399) );
  XOR U428 ( .A(n468), .B(n469), .Z(n396) );
  ANDN U429 ( .A(n470), .B(n471), .Z(n469) );
  XNOR U430 ( .A(n468), .B(n472), .Z(n470) );
  XOR U431 ( .A(n406), .B(n473), .Z(n400) );
  IV U432 ( .A(n405), .Z(n473) );
  XNOR U433 ( .A(n402), .B(n467), .Z(n405) );
  AND U434 ( .A(n552), .B(n395), .Z(n467) );
  XOR U435 ( .A(n474), .B(n475), .Z(n402) );
  ANDN U436 ( .A(n476), .B(n477), .Z(n475) );
  XNOR U437 ( .A(n474), .B(n478), .Z(n476) );
  XOR U438 ( .A(n412), .B(n479), .Z(n406) );
  IV U439 ( .A(n411), .Z(n479) );
  XNOR U440 ( .A(n408), .B(n460), .Z(n411) );
  AND U441 ( .A(n736), .B(n264), .Z(n460) );
  XOR U442 ( .A(n480), .B(n481), .Z(n408) );
  ANDN U443 ( .A(n482), .B(n483), .Z(n481) );
  XNOR U444 ( .A(n480), .B(n484), .Z(n482) );
  XOR U445 ( .A(n418), .B(n485), .Z(n412) );
  IV U446 ( .A(n417), .Z(n485) );
  XNOR U447 ( .A(n414), .B(n453), .Z(n417) );
  AND U448 ( .A(n948), .B(n159), .Z(n453) );
  XOR U449 ( .A(n486), .B(n487), .Z(n414) );
  ANDN U450 ( .A(n488), .B(n489), .Z(n487) );
  XNOR U451 ( .A(n486), .B(n490), .Z(n488) );
  XOR U452 ( .A(n425), .B(n491), .Z(n418) );
  IV U453 ( .A(n424), .Z(n491) );
  XNOR U454 ( .A(n421), .B(n446), .Z(n424) );
  AND U455 ( .A(n1185), .B(n80), .Z(n446) );
  XOR U456 ( .A(n492), .B(n493), .Z(n421) );
  ANDN U457 ( .A(n494), .B(n495), .Z(n493) );
  XNOR U458 ( .A(n492), .B(n496), .Z(n494) );
  XOR U459 ( .A(n430), .B(n497), .Z(n425) );
  IV U460 ( .A(n429), .Z(n497) );
  XNOR U461 ( .A(n426), .B(n498), .Z(n429) );
  AND U462 ( .A(n42), .B(n1448), .Z(n498) );
  XOR U463 ( .A(n499), .B(n500), .Z(n426) );
  ANDN U464 ( .A(n501), .B(n502), .Z(n500) );
  XNOR U465 ( .A(n499), .B(n503), .Z(n501) );
  XNOR U466 ( .A(n504), .B(n505), .Z(n430) );
  ANDN U467 ( .A(n506), .B(n507), .Z(n505) );
  XNOR U468 ( .A(n504), .B(n508), .Z(n506) );
  XNOR U469 ( .A(n438), .B(n431), .Z(n444) );
  XOR U470 ( .A(n509), .B(n510), .Z(n431) );
  AND U471 ( .A(n511), .B(n512), .Z(n510) );
  XNOR U472 ( .A(n9), .B(n509), .Z(n512) );
  XOR U473 ( .A(n436), .B(n513), .Z(n438) );
  ANDN U474 ( .A(n1448), .B(n43), .Z(n513) );
  XOR U475 ( .A(n514), .B(n515), .Z(n436) );
  AND U476 ( .A(n516), .B(n517), .Z(n515) );
  XNOR U477 ( .A(n514), .B(n518), .Z(n517) );
  NANDN U478 ( .B(n519), .A(n520), .Z(n441) );
  NANDN U479 ( .B(n519), .A(n521), .Z(n520) );
  XNOR U480 ( .A(n9), .B(n511), .Z(n521) );
  XOR U481 ( .A(n522), .B(n518), .Z(n511) );
  XOR U482 ( .A(n451), .B(n523), .Z(n518) );
  IV U483 ( .A(n450), .Z(n523) );
  XNOR U484 ( .A(n447), .B(n524), .Z(n450) );
  XOR U485 ( .A(n525), .B(n526), .Z(n447) );
  ANDN U486 ( .A(n527), .B(n528), .Z(n526) );
  XNOR U487 ( .A(n525), .B(n529), .Z(n527) );
  XOR U488 ( .A(n458), .B(n530), .Z(n451) );
  IV U489 ( .A(n457), .Z(n530) );
  XNOR U490 ( .A(n454), .B(n531), .Z(n457) );
  XOR U491 ( .A(n532), .B(n533), .Z(n454) );
  ANDN U492 ( .A(n534), .B(n535), .Z(n533) );
  XNOR U493 ( .A(n532), .B(n536), .Z(n534) );
  XOR U494 ( .A(n465), .B(n537), .Z(n458) );
  IV U495 ( .A(n464), .Z(n537) );
  XNOR U496 ( .A(n461), .B(n538), .Z(n464) );
  XOR U497 ( .A(n539), .B(n540), .Z(n461) );
  ANDN U498 ( .A(n541), .B(n542), .Z(n540) );
  XNOR U499 ( .A(n539), .B(n543), .Z(n541) );
  XOR U500 ( .A(n472), .B(n544), .Z(n465) );
  IV U501 ( .A(n471), .Z(n544) );
  XNOR U502 ( .A(n468), .B(n545), .Z(n471) );
  XOR U503 ( .A(n546), .B(n547), .Z(n468) );
  ANDN U504 ( .A(n548), .B(n549), .Z(n547) );
  XNOR U505 ( .A(n546), .B(n550), .Z(n548) );
  XOR U506 ( .A(n478), .B(n551), .Z(n472) );
  IV U507 ( .A(n477), .Z(n551) );
  XNOR U508 ( .A(n474), .B(n552), .Z(n477) );
  XOR U509 ( .A(n553), .B(n554), .Z(n474) );
  ANDN U510 ( .A(n555), .B(n556), .Z(n554) );
  XNOR U511 ( .A(n553), .B(n557), .Z(n555) );
  XOR U512 ( .A(n484), .B(n558), .Z(n478) );
  IV U513 ( .A(n483), .Z(n558) );
  XNOR U514 ( .A(n480), .B(n545), .Z(n483) );
  AND U515 ( .A(n736), .B(n395), .Z(n545) );
  XOR U516 ( .A(n559), .B(n560), .Z(n480) );
  ANDN U517 ( .A(n561), .B(n562), .Z(n560) );
  XNOR U518 ( .A(n559), .B(n563), .Z(n561) );
  XOR U519 ( .A(n490), .B(n564), .Z(n484) );
  IV U520 ( .A(n489), .Z(n564) );
  XNOR U521 ( .A(n486), .B(n538), .Z(n489) );
  AND U522 ( .A(n948), .B(n264), .Z(n538) );
  XOR U523 ( .A(n565), .B(n566), .Z(n486) );
  ANDN U524 ( .A(n567), .B(n568), .Z(n566) );
  XNOR U525 ( .A(n565), .B(n569), .Z(n567) );
  XOR U526 ( .A(n496), .B(n570), .Z(n490) );
  IV U527 ( .A(n495), .Z(n570) );
  XNOR U528 ( .A(n492), .B(n531), .Z(n495) );
  AND U529 ( .A(n1185), .B(n159), .Z(n531) );
  XOR U530 ( .A(n571), .B(n572), .Z(n492) );
  ANDN U531 ( .A(n573), .B(n574), .Z(n572) );
  XNOR U532 ( .A(n571), .B(n575), .Z(n573) );
  XOR U533 ( .A(n503), .B(n576), .Z(n496) );
  IV U534 ( .A(n502), .Z(n576) );
  XNOR U535 ( .A(n499), .B(n524), .Z(n502) );
  AND U536 ( .A(n1448), .B(n80), .Z(n524) );
  XOR U537 ( .A(n577), .B(n578), .Z(n499) );
  ANDN U538 ( .A(n579), .B(n580), .Z(n578) );
  XNOR U539 ( .A(n577), .B(n581), .Z(n579) );
  XOR U540 ( .A(n508), .B(n582), .Z(n503) );
  IV U541 ( .A(n507), .Z(n582) );
  XNOR U542 ( .A(n504), .B(n583), .Z(n507) );
  AND U543 ( .A(n42), .B(n1737), .Z(n583) );
  XOR U544 ( .A(n584), .B(n585), .Z(n504) );
  ANDN U545 ( .A(n586), .B(n587), .Z(n585) );
  XNOR U546 ( .A(n584), .B(n588), .Z(n586) );
  XNOR U547 ( .A(n589), .B(n590), .Z(n508) );
  ANDN U548 ( .A(n591), .B(n592), .Z(n590) );
  XNOR U549 ( .A(n589), .B(n593), .Z(n591) );
  XNOR U550 ( .A(n516), .B(n509), .Z(n522) );
  XOR U551 ( .A(n594), .B(n595), .Z(n509) );
  AND U552 ( .A(n596), .B(n597), .Z(n595) );
  XNOR U553 ( .A(n9), .B(n594), .Z(n597) );
  XOR U554 ( .A(n514), .B(n598), .Z(n516) );
  ANDN U555 ( .A(n1737), .B(n43), .Z(n598) );
  XOR U556 ( .A(n599), .B(n600), .Z(n514) );
  AND U557 ( .A(n601), .B(n602), .Z(n600) );
  XNOR U558 ( .A(n599), .B(n603), .Z(n602) );
  NANDN U559 ( .B(n604), .A(n605), .Z(n519) );
  NANDN U560 ( .B(n604), .A(n606), .Z(n605) );
  XNOR U561 ( .A(n9), .B(n596), .Z(n606) );
  XOR U562 ( .A(n607), .B(n603), .Z(n596) );
  XOR U563 ( .A(n529), .B(n608), .Z(n603) );
  IV U564 ( .A(n528), .Z(n608) );
  XNOR U565 ( .A(n525), .B(n609), .Z(n528) );
  XOR U566 ( .A(n610), .B(n611), .Z(n525) );
  ANDN U567 ( .A(n612), .B(n613), .Z(n611) );
  XNOR U568 ( .A(n610), .B(n614), .Z(n612) );
  XOR U569 ( .A(n536), .B(n615), .Z(n529) );
  IV U570 ( .A(n535), .Z(n615) );
  XNOR U571 ( .A(n532), .B(n616), .Z(n535) );
  XOR U572 ( .A(n617), .B(n618), .Z(n532) );
  ANDN U573 ( .A(n619), .B(n620), .Z(n618) );
  XNOR U574 ( .A(n617), .B(n621), .Z(n619) );
  XOR U575 ( .A(n543), .B(n622), .Z(n536) );
  IV U576 ( .A(n542), .Z(n622) );
  XNOR U577 ( .A(n539), .B(n623), .Z(n542) );
  XOR U578 ( .A(n624), .B(n625), .Z(n539) );
  ANDN U579 ( .A(n626), .B(n627), .Z(n625) );
  XNOR U580 ( .A(n624), .B(n628), .Z(n626) );
  XOR U581 ( .A(n550), .B(n629), .Z(n543) );
  IV U582 ( .A(n549), .Z(n629) );
  XNOR U583 ( .A(n546), .B(n630), .Z(n549) );
  XOR U584 ( .A(n631), .B(n632), .Z(n546) );
  ANDN U585 ( .A(n633), .B(n634), .Z(n632) );
  XNOR U586 ( .A(n631), .B(n635), .Z(n633) );
  XOR U587 ( .A(n557), .B(n636), .Z(n550) );
  IV U588 ( .A(n556), .Z(n636) );
  XNOR U589 ( .A(n553), .B(n637), .Z(n556) );
  XOR U590 ( .A(n638), .B(n639), .Z(n553) );
  ANDN U591 ( .A(n640), .B(n641), .Z(n639) );
  XNOR U592 ( .A(n638), .B(n642), .Z(n640) );
  XOR U593 ( .A(n563), .B(n643), .Z(n557) );
  IV U594 ( .A(n562), .Z(n643) );
  XNOR U595 ( .A(n559), .B(n637), .Z(n562) );
  AND U596 ( .A(n736), .B(n552), .Z(n637) );
  XOR U597 ( .A(n644), .B(n645), .Z(n559) );
  ANDN U598 ( .A(n646), .B(n647), .Z(n645) );
  XNOR U599 ( .A(n644), .B(n648), .Z(n646) );
  XOR U600 ( .A(n569), .B(n649), .Z(n563) );
  IV U601 ( .A(n568), .Z(n649) );
  XNOR U602 ( .A(n565), .B(n630), .Z(n568) );
  AND U603 ( .A(n948), .B(n395), .Z(n630) );
  XOR U604 ( .A(n650), .B(n651), .Z(n565) );
  ANDN U605 ( .A(n652), .B(n653), .Z(n651) );
  XNOR U606 ( .A(n650), .B(n654), .Z(n652) );
  XOR U607 ( .A(n575), .B(n655), .Z(n569) );
  IV U608 ( .A(n574), .Z(n655) );
  XNOR U609 ( .A(n571), .B(n623), .Z(n574) );
  AND U610 ( .A(n1185), .B(n264), .Z(n623) );
  XOR U611 ( .A(n656), .B(n657), .Z(n571) );
  ANDN U612 ( .A(n658), .B(n659), .Z(n657) );
  XNOR U613 ( .A(n656), .B(n660), .Z(n658) );
  XOR U614 ( .A(n581), .B(n661), .Z(n575) );
  IV U615 ( .A(n580), .Z(n661) );
  XNOR U616 ( .A(n577), .B(n616), .Z(n580) );
  AND U617 ( .A(n1448), .B(n159), .Z(n616) );
  XOR U618 ( .A(n662), .B(n663), .Z(n577) );
  ANDN U619 ( .A(n664), .B(n665), .Z(n663) );
  XNOR U620 ( .A(n662), .B(n666), .Z(n664) );
  XOR U621 ( .A(n588), .B(n667), .Z(n581) );
  IV U622 ( .A(n587), .Z(n667) );
  XNOR U623 ( .A(n584), .B(n609), .Z(n587) );
  AND U624 ( .A(n1737), .B(n80), .Z(n609) );
  XOR U625 ( .A(n668), .B(n669), .Z(n584) );
  ANDN U626 ( .A(n670), .B(n671), .Z(n669) );
  XNOR U627 ( .A(n668), .B(n672), .Z(n670) );
  XOR U628 ( .A(n593), .B(n673), .Z(n588) );
  IV U629 ( .A(n592), .Z(n673) );
  XNOR U630 ( .A(n589), .B(n674), .Z(n592) );
  AND U631 ( .A(n42), .B(n2053), .Z(n674) );
  XOR U632 ( .A(n675), .B(n676), .Z(n589) );
  ANDN U633 ( .A(n677), .B(n678), .Z(n676) );
  XNOR U634 ( .A(n675), .B(n679), .Z(n677) );
  XNOR U635 ( .A(n680), .B(n681), .Z(n593) );
  ANDN U636 ( .A(n682), .B(n683), .Z(n681) );
  XNOR U637 ( .A(n680), .B(n684), .Z(n682) );
  XNOR U638 ( .A(n601), .B(n594), .Z(n607) );
  XOR U639 ( .A(n685), .B(n686), .Z(n594) );
  AND U640 ( .A(n687), .B(n688), .Z(n686) );
  XNOR U641 ( .A(n9), .B(n685), .Z(n688) );
  XOR U642 ( .A(n599), .B(n689), .Z(n601) );
  ANDN U643 ( .A(n2053), .B(n43), .Z(n689) );
  XOR U644 ( .A(n690), .B(n691), .Z(n599) );
  AND U645 ( .A(n692), .B(n693), .Z(n691) );
  XNOR U646 ( .A(n690), .B(n694), .Z(n693) );
  NAND U647 ( .A(n695), .B(n696), .Z(n604) );
  NAND U648 ( .A(n697), .B(n696), .Z(n695) );
  XOR U649 ( .A(n698), .B(n687), .Z(n697) );
  XOR U650 ( .A(n699), .B(n694), .Z(n687) );
  XOR U651 ( .A(n614), .B(n700), .Z(n694) );
  IV U652 ( .A(n613), .Z(n700) );
  XNOR U653 ( .A(n610), .B(n701), .Z(n613) );
  XOR U654 ( .A(n702), .B(n703), .Z(n610) );
  ANDN U655 ( .A(n704), .B(n705), .Z(n703) );
  XNOR U656 ( .A(n702), .B(n706), .Z(n704) );
  XOR U657 ( .A(n621), .B(n707), .Z(n614) );
  IV U658 ( .A(n620), .Z(n707) );
  XNOR U659 ( .A(n617), .B(n708), .Z(n620) );
  XOR U660 ( .A(n709), .B(n710), .Z(n617) );
  ANDN U661 ( .A(n711), .B(n712), .Z(n710) );
  XNOR U662 ( .A(n709), .B(n713), .Z(n711) );
  XOR U663 ( .A(n628), .B(n714), .Z(n621) );
  IV U664 ( .A(n627), .Z(n714) );
  XNOR U665 ( .A(n624), .B(n715), .Z(n627) );
  XOR U666 ( .A(n716), .B(n717), .Z(n624) );
  ANDN U667 ( .A(n718), .B(n719), .Z(n717) );
  XNOR U668 ( .A(n716), .B(n720), .Z(n718) );
  XOR U669 ( .A(n635), .B(n721), .Z(n628) );
  IV U670 ( .A(n634), .Z(n721) );
  XNOR U671 ( .A(n631), .B(n722), .Z(n634) );
  XOR U672 ( .A(n723), .B(n724), .Z(n631) );
  ANDN U673 ( .A(n725), .B(n726), .Z(n724) );
  XNOR U674 ( .A(n723), .B(n727), .Z(n725) );
  XOR U675 ( .A(n642), .B(n728), .Z(n635) );
  IV U676 ( .A(n641), .Z(n728) );
  XNOR U677 ( .A(n638), .B(n729), .Z(n641) );
  XOR U678 ( .A(n730), .B(n731), .Z(n638) );
  ANDN U679 ( .A(n732), .B(n733), .Z(n731) );
  XNOR U680 ( .A(n730), .B(n734), .Z(n732) );
  XOR U681 ( .A(n648), .B(n735), .Z(n642) );
  IV U682 ( .A(n647), .Z(n735) );
  XNOR U683 ( .A(n644), .B(n736), .Z(n647) );
  XOR U684 ( .A(n737), .B(n738), .Z(n644) );
  ANDN U685 ( .A(n739), .B(n740), .Z(n738) );
  XNOR U686 ( .A(n737), .B(n741), .Z(n739) );
  XOR U687 ( .A(n654), .B(n742), .Z(n648) );
  IV U688 ( .A(n653), .Z(n742) );
  XNOR U689 ( .A(n650), .B(n729), .Z(n653) );
  AND U690 ( .A(n948), .B(n552), .Z(n729) );
  XOR U691 ( .A(n743), .B(n744), .Z(n650) );
  ANDN U692 ( .A(n745), .B(n746), .Z(n744) );
  XNOR U693 ( .A(n743), .B(n747), .Z(n745) );
  XOR U694 ( .A(n660), .B(n748), .Z(n654) );
  IV U695 ( .A(n659), .Z(n748) );
  XNOR U696 ( .A(n656), .B(n722), .Z(n659) );
  AND U697 ( .A(n1185), .B(n395), .Z(n722) );
  XOR U698 ( .A(n749), .B(n750), .Z(n656) );
  ANDN U699 ( .A(n751), .B(n752), .Z(n750) );
  XNOR U700 ( .A(n749), .B(n753), .Z(n751) );
  XOR U701 ( .A(n666), .B(n754), .Z(n660) );
  IV U702 ( .A(n665), .Z(n754) );
  XNOR U703 ( .A(n662), .B(n715), .Z(n665) );
  AND U704 ( .A(n1448), .B(n264), .Z(n715) );
  XOR U705 ( .A(n755), .B(n756), .Z(n662) );
  ANDN U706 ( .A(n757), .B(n758), .Z(n756) );
  XNOR U707 ( .A(n755), .B(n759), .Z(n757) );
  XOR U708 ( .A(n672), .B(n760), .Z(n666) );
  IV U709 ( .A(n671), .Z(n760) );
  XNOR U710 ( .A(n668), .B(n708), .Z(n671) );
  AND U711 ( .A(n1737), .B(n159), .Z(n708) );
  XOR U712 ( .A(n761), .B(n762), .Z(n668) );
  ANDN U713 ( .A(n763), .B(n764), .Z(n762) );
  XNOR U714 ( .A(n761), .B(n765), .Z(n763) );
  XOR U715 ( .A(n679), .B(n766), .Z(n672) );
  IV U716 ( .A(n678), .Z(n766) );
  XNOR U717 ( .A(n675), .B(n701), .Z(n678) );
  AND U718 ( .A(n2053), .B(n80), .Z(n701) );
  XOR U719 ( .A(n767), .B(n768), .Z(n675) );
  ANDN U720 ( .A(n769), .B(n770), .Z(n768) );
  XNOR U721 ( .A(n767), .B(n771), .Z(n769) );
  XOR U722 ( .A(n684), .B(n772), .Z(n679) );
  IV U723 ( .A(n683), .Z(n772) );
  XNOR U724 ( .A(n680), .B(n773), .Z(n683) );
  AND U725 ( .A(n42), .B(n2396), .Z(n773) );
  XOR U726 ( .A(n774), .B(n775), .Z(n680) );
  ANDN U727 ( .A(n776), .B(n777), .Z(n775) );
  XNOR U728 ( .A(n774), .B(n778), .Z(n776) );
  XNOR U729 ( .A(n779), .B(n780), .Z(n684) );
  ANDN U730 ( .A(n781), .B(n782), .Z(n780) );
  XNOR U731 ( .A(n779), .B(n783), .Z(n781) );
  XNOR U732 ( .A(n692), .B(n685), .Z(n699) );
  XOR U733 ( .A(n784), .B(n785), .Z(n685) );
  AND U734 ( .A(n786), .B(n787), .Z(n785) );
  XNOR U735 ( .A(n9), .B(n784), .Z(n787) );
  XOR U736 ( .A(n690), .B(n788), .Z(n692) );
  ANDN U737 ( .A(n2396), .B(n43), .Z(n788) );
  XOR U738 ( .A(n789), .B(n790), .Z(n690) );
  AND U739 ( .A(n791), .B(n792), .Z(n790) );
  XNOR U740 ( .A(n789), .B(n793), .Z(n792) );
  XNOR U741 ( .A(n794), .B(n696), .Z(n698) );
  AND U742 ( .A(n795), .B(n796), .Z(n696) );
  NAND U743 ( .A(n797), .B(n796), .Z(n795) );
  XOR U744 ( .A(n798), .B(n786), .Z(n797) );
  XOR U745 ( .A(n799), .B(n793), .Z(n786) );
  XOR U746 ( .A(n706), .B(n800), .Z(n793) );
  IV U747 ( .A(n705), .Z(n800) );
  XNOR U748 ( .A(n702), .B(n801), .Z(n705) );
  XOR U749 ( .A(n802), .B(n803), .Z(n702) );
  ANDN U750 ( .A(n804), .B(n805), .Z(n803) );
  XNOR U751 ( .A(n802), .B(n806), .Z(n804) );
  XOR U752 ( .A(n713), .B(n807), .Z(n706) );
  IV U753 ( .A(n712), .Z(n807) );
  XNOR U754 ( .A(n709), .B(n808), .Z(n712) );
  XOR U755 ( .A(n809), .B(n810), .Z(n709) );
  ANDN U756 ( .A(n811), .B(n812), .Z(n810) );
  XNOR U757 ( .A(n809), .B(n813), .Z(n811) );
  XOR U758 ( .A(n720), .B(n814), .Z(n713) );
  IV U759 ( .A(n719), .Z(n814) );
  XNOR U760 ( .A(n716), .B(n815), .Z(n719) );
  XOR U761 ( .A(n816), .B(n817), .Z(n716) );
  ANDN U762 ( .A(n818), .B(n819), .Z(n817) );
  XNOR U763 ( .A(n816), .B(n820), .Z(n818) );
  XOR U764 ( .A(n727), .B(n821), .Z(n720) );
  IV U765 ( .A(n726), .Z(n821) );
  XNOR U766 ( .A(n723), .B(n822), .Z(n726) );
  XOR U767 ( .A(n823), .B(n824), .Z(n723) );
  ANDN U768 ( .A(n825), .B(n826), .Z(n824) );
  XNOR U769 ( .A(n823), .B(n827), .Z(n825) );
  XOR U770 ( .A(n734), .B(n828), .Z(n727) );
  IV U771 ( .A(n733), .Z(n828) );
  XNOR U772 ( .A(n730), .B(n829), .Z(n733) );
  XOR U773 ( .A(n830), .B(n831), .Z(n730) );
  ANDN U774 ( .A(n832), .B(n833), .Z(n831) );
  XNOR U775 ( .A(n830), .B(n834), .Z(n832) );
  XOR U776 ( .A(n741), .B(n835), .Z(n734) );
  IV U777 ( .A(n740), .Z(n835) );
  XNOR U778 ( .A(n737), .B(n836), .Z(n740) );
  XOR U779 ( .A(n837), .B(n838), .Z(n737) );
  ANDN U780 ( .A(n839), .B(n840), .Z(n838) );
  XNOR U781 ( .A(n837), .B(n841), .Z(n839) );
  XOR U782 ( .A(n747), .B(n842), .Z(n741) );
  IV U783 ( .A(n746), .Z(n842) );
  XNOR U784 ( .A(n743), .B(n836), .Z(n746) );
  AND U785 ( .A(n948), .B(n736), .Z(n836) );
  XOR U786 ( .A(n843), .B(n844), .Z(n743) );
  ANDN U787 ( .A(n845), .B(n846), .Z(n844) );
  XNOR U788 ( .A(n843), .B(n847), .Z(n845) );
  XOR U789 ( .A(n753), .B(n848), .Z(n747) );
  IV U790 ( .A(n752), .Z(n848) );
  XNOR U791 ( .A(n749), .B(n829), .Z(n752) );
  AND U792 ( .A(n1185), .B(n552), .Z(n829) );
  XOR U793 ( .A(n849), .B(n850), .Z(n749) );
  ANDN U794 ( .A(n851), .B(n852), .Z(n850) );
  XNOR U795 ( .A(n849), .B(n853), .Z(n851) );
  XOR U796 ( .A(n759), .B(n854), .Z(n753) );
  IV U797 ( .A(n758), .Z(n854) );
  XNOR U798 ( .A(n755), .B(n822), .Z(n758) );
  AND U799 ( .A(n1448), .B(n395), .Z(n822) );
  XOR U800 ( .A(n855), .B(n856), .Z(n755) );
  ANDN U801 ( .A(n857), .B(n858), .Z(n856) );
  XNOR U802 ( .A(n855), .B(n859), .Z(n857) );
  XOR U803 ( .A(n765), .B(n860), .Z(n759) );
  IV U804 ( .A(n764), .Z(n860) );
  XNOR U805 ( .A(n761), .B(n815), .Z(n764) );
  AND U806 ( .A(n1737), .B(n264), .Z(n815) );
  XOR U807 ( .A(n861), .B(n862), .Z(n761) );
  ANDN U808 ( .A(n863), .B(n864), .Z(n862) );
  XNOR U809 ( .A(n861), .B(n865), .Z(n863) );
  XOR U810 ( .A(n771), .B(n866), .Z(n765) );
  IV U811 ( .A(n770), .Z(n866) );
  XNOR U812 ( .A(n767), .B(n808), .Z(n770) );
  AND U813 ( .A(n2053), .B(n159), .Z(n808) );
  XOR U814 ( .A(n867), .B(n868), .Z(n767) );
  ANDN U815 ( .A(n869), .B(n870), .Z(n868) );
  XNOR U816 ( .A(n867), .B(n871), .Z(n869) );
  XOR U817 ( .A(n778), .B(n872), .Z(n771) );
  IV U818 ( .A(n777), .Z(n872) );
  XNOR U819 ( .A(n774), .B(n801), .Z(n777) );
  AND U820 ( .A(n2396), .B(n80), .Z(n801) );
  XOR U821 ( .A(n873), .B(n874), .Z(n774) );
  ANDN U822 ( .A(n875), .B(n876), .Z(n874) );
  XNOR U823 ( .A(n873), .B(n877), .Z(n875) );
  XOR U824 ( .A(n783), .B(n878), .Z(n778) );
  IV U825 ( .A(n782), .Z(n878) );
  XNOR U826 ( .A(n779), .B(n879), .Z(n782) );
  AND U827 ( .A(n42), .B(n2765), .Z(n879) );
  XOR U828 ( .A(n880), .B(n881), .Z(n779) );
  ANDN U829 ( .A(n882), .B(n883), .Z(n881) );
  XNOR U830 ( .A(n880), .B(n884), .Z(n882) );
  XNOR U831 ( .A(n885), .B(n886), .Z(n783) );
  ANDN U832 ( .A(n887), .B(n888), .Z(n886) );
  XNOR U833 ( .A(n885), .B(n889), .Z(n887) );
  XNOR U834 ( .A(n791), .B(n784), .Z(n799) );
  XOR U835 ( .A(n890), .B(n891), .Z(n784) );
  AND U836 ( .A(n892), .B(n893), .Z(n891) );
  XNOR U837 ( .A(n9), .B(n890), .Z(n893) );
  XOR U838 ( .A(n789), .B(n894), .Z(n791) );
  ANDN U839 ( .A(n2765), .B(n43), .Z(n894) );
  XOR U840 ( .A(n895), .B(n896), .Z(n789) );
  AND U841 ( .A(n897), .B(n898), .Z(n896) );
  XNOR U842 ( .A(n895), .B(n899), .Z(n898) );
  XNOR U843 ( .A(n794), .B(n796), .Z(n798) );
  AND U844 ( .A(n900), .B(n901), .Z(n796) );
  NAND U845 ( .A(n902), .B(n901), .Z(n900) );
  XOR U846 ( .A(n903), .B(n892), .Z(n902) );
  XOR U847 ( .A(n904), .B(n899), .Z(n892) );
  XOR U848 ( .A(n806), .B(n905), .Z(n899) );
  IV U849 ( .A(n805), .Z(n905) );
  XNOR U850 ( .A(n802), .B(n906), .Z(n805) );
  XOR U851 ( .A(n907), .B(n908), .Z(n802) );
  ANDN U852 ( .A(n909), .B(n910), .Z(n908) );
  XNOR U853 ( .A(n907), .B(n911), .Z(n909) );
  XOR U854 ( .A(n813), .B(n912), .Z(n806) );
  IV U855 ( .A(n812), .Z(n912) );
  XNOR U856 ( .A(n809), .B(n913), .Z(n812) );
  XOR U857 ( .A(n914), .B(n915), .Z(n809) );
  ANDN U858 ( .A(n916), .B(n917), .Z(n915) );
  XNOR U859 ( .A(n914), .B(n918), .Z(n916) );
  XOR U860 ( .A(n820), .B(n919), .Z(n813) );
  IV U861 ( .A(n819), .Z(n919) );
  XNOR U862 ( .A(n816), .B(n920), .Z(n819) );
  XOR U863 ( .A(n921), .B(n922), .Z(n816) );
  ANDN U864 ( .A(n923), .B(n924), .Z(n922) );
  XNOR U865 ( .A(n921), .B(n925), .Z(n923) );
  XOR U866 ( .A(n827), .B(n926), .Z(n820) );
  IV U867 ( .A(n826), .Z(n926) );
  XNOR U868 ( .A(n823), .B(n927), .Z(n826) );
  XOR U869 ( .A(n928), .B(n929), .Z(n823) );
  ANDN U870 ( .A(n930), .B(n931), .Z(n929) );
  XNOR U871 ( .A(n928), .B(n932), .Z(n930) );
  XOR U872 ( .A(n834), .B(n933), .Z(n827) );
  IV U873 ( .A(n833), .Z(n933) );
  XNOR U874 ( .A(n830), .B(n934), .Z(n833) );
  XOR U875 ( .A(n935), .B(n936), .Z(n830) );
  ANDN U876 ( .A(n937), .B(n938), .Z(n936) );
  XNOR U877 ( .A(n935), .B(n939), .Z(n937) );
  XOR U878 ( .A(n841), .B(n940), .Z(n834) );
  IV U879 ( .A(n840), .Z(n940) );
  XNOR U880 ( .A(n837), .B(n941), .Z(n840) );
  XOR U881 ( .A(n942), .B(n943), .Z(n837) );
  ANDN U882 ( .A(n944), .B(n945), .Z(n943) );
  XNOR U883 ( .A(n942), .B(n946), .Z(n944) );
  XOR U884 ( .A(n847), .B(n947), .Z(n841) );
  IV U885 ( .A(n846), .Z(n947) );
  XNOR U886 ( .A(n843), .B(n948), .Z(n846) );
  XOR U887 ( .A(n949), .B(n950), .Z(n843) );
  ANDN U888 ( .A(n951), .B(n952), .Z(n950) );
  XNOR U889 ( .A(n949), .B(n953), .Z(n951) );
  XOR U890 ( .A(n853), .B(n954), .Z(n847) );
  IV U891 ( .A(n852), .Z(n954) );
  XNOR U892 ( .A(n849), .B(n941), .Z(n852) );
  AND U893 ( .A(n1185), .B(n736), .Z(n941) );
  XOR U894 ( .A(n955), .B(n956), .Z(n849) );
  ANDN U895 ( .A(n957), .B(n958), .Z(n956) );
  XNOR U896 ( .A(n955), .B(n959), .Z(n957) );
  XOR U897 ( .A(n859), .B(n960), .Z(n853) );
  IV U898 ( .A(n858), .Z(n960) );
  XNOR U899 ( .A(n855), .B(n934), .Z(n858) );
  AND U900 ( .A(n1448), .B(n552), .Z(n934) );
  XOR U901 ( .A(n961), .B(n962), .Z(n855) );
  ANDN U902 ( .A(n963), .B(n964), .Z(n962) );
  XNOR U903 ( .A(n961), .B(n965), .Z(n963) );
  XOR U904 ( .A(n865), .B(n966), .Z(n859) );
  IV U905 ( .A(n864), .Z(n966) );
  XNOR U906 ( .A(n861), .B(n927), .Z(n864) );
  AND U907 ( .A(n1737), .B(n395), .Z(n927) );
  XOR U908 ( .A(n967), .B(n968), .Z(n861) );
  ANDN U909 ( .A(n969), .B(n970), .Z(n968) );
  XNOR U910 ( .A(n967), .B(n971), .Z(n969) );
  XOR U911 ( .A(n871), .B(n972), .Z(n865) );
  IV U912 ( .A(n870), .Z(n972) );
  XNOR U913 ( .A(n867), .B(n920), .Z(n870) );
  AND U914 ( .A(n2053), .B(n264), .Z(n920) );
  XOR U915 ( .A(n973), .B(n974), .Z(n867) );
  ANDN U916 ( .A(n975), .B(n976), .Z(n974) );
  XNOR U917 ( .A(n973), .B(n977), .Z(n975) );
  XOR U918 ( .A(n877), .B(n978), .Z(n871) );
  IV U919 ( .A(n876), .Z(n978) );
  XNOR U920 ( .A(n873), .B(n913), .Z(n876) );
  AND U921 ( .A(n2396), .B(n159), .Z(n913) );
  XOR U922 ( .A(n979), .B(n980), .Z(n873) );
  ANDN U923 ( .A(n981), .B(n982), .Z(n980) );
  XNOR U924 ( .A(n979), .B(n983), .Z(n981) );
  XOR U925 ( .A(n884), .B(n984), .Z(n877) );
  IV U926 ( .A(n883), .Z(n984) );
  XNOR U927 ( .A(n880), .B(n906), .Z(n883) );
  AND U928 ( .A(n2765), .B(n80), .Z(n906) );
  XOR U929 ( .A(n985), .B(n986), .Z(n880) );
  ANDN U930 ( .A(n987), .B(n988), .Z(n986) );
  XNOR U931 ( .A(n985), .B(n989), .Z(n987) );
  XOR U932 ( .A(n889), .B(n990), .Z(n884) );
  IV U933 ( .A(n888), .Z(n990) );
  XNOR U934 ( .A(n885), .B(n991), .Z(n888) );
  AND U935 ( .A(n42), .B(n3166), .Z(n991) );
  XOR U936 ( .A(n992), .B(n993), .Z(n885) );
  ANDN U937 ( .A(n994), .B(n995), .Z(n993) );
  XNOR U938 ( .A(n992), .B(n996), .Z(n994) );
  XNOR U939 ( .A(n997), .B(n998), .Z(n889) );
  ANDN U940 ( .A(n999), .B(n1000), .Z(n998) );
  XNOR U941 ( .A(n997), .B(n1001), .Z(n999) );
  XNOR U942 ( .A(n897), .B(n890), .Z(n904) );
  XOR U943 ( .A(n1002), .B(n1003), .Z(n890) );
  AND U944 ( .A(n1004), .B(n1005), .Z(n1003) );
  XNOR U945 ( .A(n9), .B(n1002), .Z(n1005) );
  XOR U946 ( .A(n895), .B(n1006), .Z(n897) );
  ANDN U947 ( .A(n3166), .B(n43), .Z(n1006) );
  XOR U948 ( .A(n1007), .B(n1008), .Z(n895) );
  AND U949 ( .A(n1009), .B(n1010), .Z(n1008) );
  XNOR U950 ( .A(n1007), .B(n1011), .Z(n1010) );
  XNOR U951 ( .A(n794), .B(n901), .Z(n903) );
  AND U952 ( .A(n1012), .B(n1013), .Z(n901) );
  NAND U953 ( .A(n1014), .B(n1013), .Z(n1012) );
  XOR U954 ( .A(n1015), .B(n1004), .Z(n1014) );
  XOR U955 ( .A(n1016), .B(n1011), .Z(n1004) );
  XOR U956 ( .A(n911), .B(n1017), .Z(n1011) );
  IV U957 ( .A(n910), .Z(n1017) );
  XNOR U958 ( .A(n907), .B(n1018), .Z(n910) );
  XOR U959 ( .A(n1019), .B(n1020), .Z(n907) );
  ANDN U960 ( .A(n1021), .B(n1022), .Z(n1020) );
  XNOR U961 ( .A(n1019), .B(n1023), .Z(n1021) );
  XOR U962 ( .A(n918), .B(n1024), .Z(n911) );
  IV U963 ( .A(n917), .Z(n1024) );
  XNOR U964 ( .A(n914), .B(n1025), .Z(n917) );
  XOR U965 ( .A(n1026), .B(n1027), .Z(n914) );
  ANDN U966 ( .A(n1028), .B(n1029), .Z(n1027) );
  XNOR U967 ( .A(n1026), .B(n1030), .Z(n1028) );
  XOR U968 ( .A(n925), .B(n1031), .Z(n918) );
  IV U969 ( .A(n924), .Z(n1031) );
  XNOR U970 ( .A(n921), .B(n1032), .Z(n924) );
  XOR U971 ( .A(n1033), .B(n1034), .Z(n921) );
  ANDN U972 ( .A(n1035), .B(n1036), .Z(n1034) );
  XNOR U973 ( .A(n1033), .B(n1037), .Z(n1035) );
  XOR U974 ( .A(n932), .B(n1038), .Z(n925) );
  IV U975 ( .A(n931), .Z(n1038) );
  XNOR U976 ( .A(n928), .B(n1039), .Z(n931) );
  XOR U977 ( .A(n1040), .B(n1041), .Z(n928) );
  ANDN U978 ( .A(n1042), .B(n1043), .Z(n1041) );
  XNOR U979 ( .A(n1040), .B(n1044), .Z(n1042) );
  XOR U980 ( .A(n939), .B(n1045), .Z(n932) );
  IV U981 ( .A(n938), .Z(n1045) );
  XNOR U982 ( .A(n935), .B(n1046), .Z(n938) );
  XOR U983 ( .A(n1047), .B(n1048), .Z(n935) );
  ANDN U984 ( .A(n1049), .B(n1050), .Z(n1048) );
  XNOR U985 ( .A(n1047), .B(n1051), .Z(n1049) );
  XOR U986 ( .A(n946), .B(n1052), .Z(n939) );
  IV U987 ( .A(n945), .Z(n1052) );
  XNOR U988 ( .A(n942), .B(n1053), .Z(n945) );
  XOR U989 ( .A(n1054), .B(n1055), .Z(n942) );
  ANDN U990 ( .A(n1056), .B(n1057), .Z(n1055) );
  XNOR U991 ( .A(n1054), .B(n1058), .Z(n1056) );
  XOR U992 ( .A(n953), .B(n1059), .Z(n946) );
  IV U993 ( .A(n952), .Z(n1059) );
  XNOR U994 ( .A(n949), .B(n1060), .Z(n952) );
  XOR U995 ( .A(n1061), .B(n1062), .Z(n949) );
  ANDN U996 ( .A(n1063), .B(n1064), .Z(n1062) );
  XNOR U997 ( .A(n1061), .B(n1065), .Z(n1063) );
  XOR U998 ( .A(n959), .B(n1066), .Z(n953) );
  IV U999 ( .A(n958), .Z(n1066) );
  XNOR U1000 ( .A(n955), .B(n1060), .Z(n958) );
  AND U1001 ( .A(n1185), .B(n948), .Z(n1060) );
  XOR U1002 ( .A(n1067), .B(n1068), .Z(n955) );
  ANDN U1003 ( .A(n1069), .B(n1070), .Z(n1068) );
  XNOR U1004 ( .A(n1067), .B(n1071), .Z(n1069) );
  XOR U1005 ( .A(n965), .B(n1072), .Z(n959) );
  IV U1006 ( .A(n964), .Z(n1072) );
  XNOR U1007 ( .A(n961), .B(n1053), .Z(n964) );
  AND U1008 ( .A(n1448), .B(n736), .Z(n1053) );
  XOR U1009 ( .A(n1073), .B(n1074), .Z(n961) );
  ANDN U1010 ( .A(n1075), .B(n1076), .Z(n1074) );
  XNOR U1011 ( .A(n1073), .B(n1077), .Z(n1075) );
  XOR U1012 ( .A(n971), .B(n1078), .Z(n965) );
  IV U1013 ( .A(n970), .Z(n1078) );
  XNOR U1014 ( .A(n967), .B(n1046), .Z(n970) );
  AND U1015 ( .A(n1737), .B(n552), .Z(n1046) );
  XOR U1016 ( .A(n1079), .B(n1080), .Z(n967) );
  ANDN U1017 ( .A(n1081), .B(n1082), .Z(n1080) );
  XNOR U1018 ( .A(n1079), .B(n1083), .Z(n1081) );
  XOR U1019 ( .A(n977), .B(n1084), .Z(n971) );
  IV U1020 ( .A(n976), .Z(n1084) );
  XNOR U1021 ( .A(n973), .B(n1039), .Z(n976) );
  AND U1022 ( .A(n2053), .B(n395), .Z(n1039) );
  XOR U1023 ( .A(n1085), .B(n1086), .Z(n973) );
  ANDN U1024 ( .A(n1087), .B(n1088), .Z(n1086) );
  XNOR U1025 ( .A(n1085), .B(n1089), .Z(n1087) );
  XOR U1026 ( .A(n983), .B(n1090), .Z(n977) );
  IV U1027 ( .A(n982), .Z(n1090) );
  XNOR U1028 ( .A(n979), .B(n1032), .Z(n982) );
  AND U1029 ( .A(n2396), .B(n264), .Z(n1032) );
  XOR U1030 ( .A(n1091), .B(n1092), .Z(n979) );
  ANDN U1031 ( .A(n1093), .B(n1094), .Z(n1092) );
  XNOR U1032 ( .A(n1091), .B(n1095), .Z(n1093) );
  XOR U1033 ( .A(n989), .B(n1096), .Z(n983) );
  IV U1034 ( .A(n988), .Z(n1096) );
  XNOR U1035 ( .A(n985), .B(n1025), .Z(n988) );
  AND U1036 ( .A(n2765), .B(n159), .Z(n1025) );
  XOR U1037 ( .A(n1097), .B(n1098), .Z(n985) );
  ANDN U1038 ( .A(n1099), .B(n1100), .Z(n1098) );
  XNOR U1039 ( .A(n1097), .B(n1101), .Z(n1099) );
  XOR U1040 ( .A(n996), .B(n1102), .Z(n989) );
  IV U1041 ( .A(n995), .Z(n1102) );
  XNOR U1042 ( .A(n992), .B(n1018), .Z(n995) );
  AND U1043 ( .A(n3166), .B(n80), .Z(n1018) );
  XOR U1044 ( .A(n1103), .B(n1104), .Z(n992) );
  ANDN U1045 ( .A(n1105), .B(n1106), .Z(n1104) );
  XNOR U1046 ( .A(n1103), .B(n1107), .Z(n1105) );
  XOR U1047 ( .A(n1001), .B(n1108), .Z(n996) );
  IV U1048 ( .A(n1000), .Z(n1108) );
  XNOR U1049 ( .A(n997), .B(n1109), .Z(n1000) );
  AND U1050 ( .A(n42), .B(n3593), .Z(n1109) );
  XOR U1051 ( .A(n1110), .B(n1111), .Z(n997) );
  ANDN U1052 ( .A(n1112), .B(n1113), .Z(n1111) );
  XNOR U1053 ( .A(n1110), .B(n1114), .Z(n1112) );
  XNOR U1054 ( .A(n1115), .B(n1116), .Z(n1001) );
  ANDN U1055 ( .A(n1117), .B(n1118), .Z(n1116) );
  XNOR U1056 ( .A(n1115), .B(n1119), .Z(n1117) );
  XNOR U1057 ( .A(n1009), .B(n1002), .Z(n1016) );
  XOR U1058 ( .A(n1120), .B(n1121), .Z(n1002) );
  AND U1059 ( .A(n1122), .B(n1123), .Z(n1121) );
  XNOR U1060 ( .A(n9), .B(n1120), .Z(n1123) );
  XOR U1061 ( .A(n1007), .B(n1124), .Z(n1009) );
  ANDN U1062 ( .A(n3593), .B(n43), .Z(n1124) );
  XOR U1063 ( .A(n1125), .B(n1126), .Z(n1007) );
  AND U1064 ( .A(n1127), .B(n1128), .Z(n1126) );
  XNOR U1065 ( .A(n1125), .B(n1129), .Z(n1128) );
  XNOR U1066 ( .A(n794), .B(n1013), .Z(n1015) );
  AND U1067 ( .A(n1130), .B(n1131), .Z(n1013) );
  NAND U1068 ( .A(n1132), .B(n1131), .Z(n1130) );
  XOR U1069 ( .A(n1133), .B(n1122), .Z(n1132) );
  XOR U1070 ( .A(n1134), .B(n1129), .Z(n1122) );
  XOR U1071 ( .A(n1023), .B(n1135), .Z(n1129) );
  IV U1072 ( .A(n1022), .Z(n1135) );
  XNOR U1073 ( .A(n1019), .B(n1136), .Z(n1022) );
  XOR U1074 ( .A(n1137), .B(n1138), .Z(n1019) );
  ANDN U1075 ( .A(n1139), .B(n1140), .Z(n1138) );
  XNOR U1076 ( .A(n1137), .B(n1141), .Z(n1139) );
  XOR U1077 ( .A(n1030), .B(n1142), .Z(n1023) );
  IV U1078 ( .A(n1029), .Z(n1142) );
  XNOR U1079 ( .A(n1026), .B(n1143), .Z(n1029) );
  XOR U1080 ( .A(n1144), .B(n1145), .Z(n1026) );
  ANDN U1081 ( .A(n1146), .B(n1147), .Z(n1145) );
  XNOR U1082 ( .A(n1144), .B(n1148), .Z(n1146) );
  XOR U1083 ( .A(n1037), .B(n1149), .Z(n1030) );
  IV U1084 ( .A(n1036), .Z(n1149) );
  XNOR U1085 ( .A(n1033), .B(n1150), .Z(n1036) );
  XOR U1086 ( .A(n1151), .B(n1152), .Z(n1033) );
  ANDN U1087 ( .A(n1153), .B(n1154), .Z(n1152) );
  XNOR U1088 ( .A(n1151), .B(n1155), .Z(n1153) );
  XOR U1089 ( .A(n1044), .B(n1156), .Z(n1037) );
  IV U1090 ( .A(n1043), .Z(n1156) );
  XNOR U1091 ( .A(n1040), .B(n1157), .Z(n1043) );
  XOR U1092 ( .A(n1158), .B(n1159), .Z(n1040) );
  ANDN U1093 ( .A(n1160), .B(n1161), .Z(n1159) );
  XNOR U1094 ( .A(n1158), .B(n1162), .Z(n1160) );
  XOR U1095 ( .A(n1051), .B(n1163), .Z(n1044) );
  IV U1096 ( .A(n1050), .Z(n1163) );
  XNOR U1097 ( .A(n1047), .B(n1164), .Z(n1050) );
  XOR U1098 ( .A(n1165), .B(n1166), .Z(n1047) );
  ANDN U1099 ( .A(n1167), .B(n1168), .Z(n1166) );
  XNOR U1100 ( .A(n1165), .B(n1169), .Z(n1167) );
  XOR U1101 ( .A(n1058), .B(n1170), .Z(n1051) );
  IV U1102 ( .A(n1057), .Z(n1170) );
  XNOR U1103 ( .A(n1054), .B(n1171), .Z(n1057) );
  XOR U1104 ( .A(n1172), .B(n1173), .Z(n1054) );
  ANDN U1105 ( .A(n1174), .B(n1175), .Z(n1173) );
  XNOR U1106 ( .A(n1172), .B(n1176), .Z(n1174) );
  XOR U1107 ( .A(n1065), .B(n1177), .Z(n1058) );
  IV U1108 ( .A(n1064), .Z(n1177) );
  XNOR U1109 ( .A(n1061), .B(n1178), .Z(n1064) );
  XOR U1110 ( .A(n1179), .B(n1180), .Z(n1061) );
  ANDN U1111 ( .A(n1181), .B(n1182), .Z(n1180) );
  XNOR U1112 ( .A(n1179), .B(n1183), .Z(n1181) );
  XOR U1113 ( .A(n1071), .B(n1184), .Z(n1065) );
  IV U1114 ( .A(n1070), .Z(n1184) );
  XNOR U1115 ( .A(n1067), .B(n1185), .Z(n1070) );
  XOR U1116 ( .A(n1186), .B(n1187), .Z(n1067) );
  ANDN U1117 ( .A(n1188), .B(n1189), .Z(n1187) );
  XNOR U1118 ( .A(n1186), .B(n1190), .Z(n1188) );
  XOR U1119 ( .A(n1077), .B(n1191), .Z(n1071) );
  IV U1120 ( .A(n1076), .Z(n1191) );
  XNOR U1121 ( .A(n1073), .B(n1178), .Z(n1076) );
  AND U1122 ( .A(n1448), .B(n948), .Z(n1178) );
  XOR U1123 ( .A(n1192), .B(n1193), .Z(n1073) );
  ANDN U1124 ( .A(n1194), .B(n1195), .Z(n1193) );
  XNOR U1125 ( .A(n1192), .B(n1196), .Z(n1194) );
  XOR U1126 ( .A(n1083), .B(n1197), .Z(n1077) );
  IV U1127 ( .A(n1082), .Z(n1197) );
  XNOR U1128 ( .A(n1079), .B(n1171), .Z(n1082) );
  AND U1129 ( .A(n1737), .B(n736), .Z(n1171) );
  XOR U1130 ( .A(n1198), .B(n1199), .Z(n1079) );
  ANDN U1131 ( .A(n1200), .B(n1201), .Z(n1199) );
  XNOR U1132 ( .A(n1198), .B(n1202), .Z(n1200) );
  XOR U1133 ( .A(n1089), .B(n1203), .Z(n1083) );
  IV U1134 ( .A(n1088), .Z(n1203) );
  XNOR U1135 ( .A(n1085), .B(n1164), .Z(n1088) );
  AND U1136 ( .A(n2053), .B(n552), .Z(n1164) );
  XOR U1137 ( .A(n1204), .B(n1205), .Z(n1085) );
  ANDN U1138 ( .A(n1206), .B(n1207), .Z(n1205) );
  XNOR U1139 ( .A(n1204), .B(n1208), .Z(n1206) );
  XOR U1140 ( .A(n1095), .B(n1209), .Z(n1089) );
  IV U1141 ( .A(n1094), .Z(n1209) );
  XNOR U1142 ( .A(n1091), .B(n1157), .Z(n1094) );
  AND U1143 ( .A(n2396), .B(n395), .Z(n1157) );
  XOR U1144 ( .A(n1210), .B(n1211), .Z(n1091) );
  ANDN U1145 ( .A(n1212), .B(n1213), .Z(n1211) );
  XNOR U1146 ( .A(n1210), .B(n1214), .Z(n1212) );
  XOR U1147 ( .A(n1101), .B(n1215), .Z(n1095) );
  IV U1148 ( .A(n1100), .Z(n1215) );
  XNOR U1149 ( .A(n1097), .B(n1150), .Z(n1100) );
  AND U1150 ( .A(n2765), .B(n264), .Z(n1150) );
  XOR U1151 ( .A(n1216), .B(n1217), .Z(n1097) );
  ANDN U1152 ( .A(n1218), .B(n1219), .Z(n1217) );
  XNOR U1153 ( .A(n1216), .B(n1220), .Z(n1218) );
  XOR U1154 ( .A(n1107), .B(n1221), .Z(n1101) );
  IV U1155 ( .A(n1106), .Z(n1221) );
  XNOR U1156 ( .A(n1103), .B(n1143), .Z(n1106) );
  AND U1157 ( .A(n3166), .B(n159), .Z(n1143) );
  XOR U1158 ( .A(n1222), .B(n1223), .Z(n1103) );
  ANDN U1159 ( .A(n1224), .B(n1225), .Z(n1223) );
  XNOR U1160 ( .A(n1222), .B(n1226), .Z(n1224) );
  XOR U1161 ( .A(n1114), .B(n1227), .Z(n1107) );
  IV U1162 ( .A(n1113), .Z(n1227) );
  XNOR U1163 ( .A(n1110), .B(n1136), .Z(n1113) );
  AND U1164 ( .A(n3593), .B(n80), .Z(n1136) );
  XOR U1165 ( .A(n1228), .B(n1229), .Z(n1110) );
  ANDN U1166 ( .A(n1230), .B(n1231), .Z(n1229) );
  XNOR U1167 ( .A(n1228), .B(n1232), .Z(n1230) );
  XOR U1168 ( .A(n1119), .B(n1233), .Z(n1114) );
  IV U1169 ( .A(n1118), .Z(n1233) );
  XNOR U1170 ( .A(n1115), .B(n1234), .Z(n1118) );
  AND U1171 ( .A(n42), .B(n4046), .Z(n1234) );
  XOR U1172 ( .A(n1235), .B(n1236), .Z(n1115) );
  ANDN U1173 ( .A(n1237), .B(n1238), .Z(n1236) );
  XNOR U1174 ( .A(n1235), .B(n1239), .Z(n1237) );
  XNOR U1175 ( .A(n1240), .B(n1241), .Z(n1119) );
  ANDN U1176 ( .A(n1242), .B(n1243), .Z(n1241) );
  XNOR U1177 ( .A(n1240), .B(n1244), .Z(n1242) );
  XNOR U1178 ( .A(n1127), .B(n1120), .Z(n1134) );
  XOR U1179 ( .A(n1245), .B(n1246), .Z(n1120) );
  AND U1180 ( .A(n1247), .B(n1248), .Z(n1246) );
  XNOR U1181 ( .A(n9), .B(n1245), .Z(n1248) );
  XOR U1182 ( .A(n1125), .B(n1249), .Z(n1127) );
  ANDN U1183 ( .A(n4046), .B(n43), .Z(n1249) );
  XOR U1184 ( .A(n1250), .B(n1251), .Z(n1125) );
  AND U1185 ( .A(n1252), .B(n1253), .Z(n1251) );
  XNOR U1186 ( .A(n1250), .B(n1254), .Z(n1253) );
  XNOR U1187 ( .A(n794), .B(n1131), .Z(n1133) );
  AND U1188 ( .A(n1255), .B(n1256), .Z(n1131) );
  NAND U1189 ( .A(n1257), .B(n1256), .Z(n1255) );
  XOR U1190 ( .A(n1258), .B(n1247), .Z(n1257) );
  XOR U1191 ( .A(n1259), .B(n1254), .Z(n1247) );
  XOR U1192 ( .A(n1141), .B(n1260), .Z(n1254) );
  IV U1193 ( .A(n1140), .Z(n1260) );
  XNOR U1194 ( .A(n1137), .B(n1261), .Z(n1140) );
  XOR U1195 ( .A(n1262), .B(n1263), .Z(n1137) );
  ANDN U1196 ( .A(n1264), .B(n1265), .Z(n1263) );
  XNOR U1197 ( .A(n1262), .B(n1266), .Z(n1264) );
  XOR U1198 ( .A(n1148), .B(n1267), .Z(n1141) );
  IV U1199 ( .A(n1147), .Z(n1267) );
  XNOR U1200 ( .A(n1144), .B(n1268), .Z(n1147) );
  XOR U1201 ( .A(n1269), .B(n1270), .Z(n1144) );
  ANDN U1202 ( .A(n1271), .B(n1272), .Z(n1270) );
  XNOR U1203 ( .A(n1269), .B(n1273), .Z(n1271) );
  XOR U1204 ( .A(n1155), .B(n1274), .Z(n1148) );
  IV U1205 ( .A(n1154), .Z(n1274) );
  XNOR U1206 ( .A(n1151), .B(n1275), .Z(n1154) );
  XOR U1207 ( .A(n1276), .B(n1277), .Z(n1151) );
  ANDN U1208 ( .A(n1278), .B(n1279), .Z(n1277) );
  XNOR U1209 ( .A(n1276), .B(n1280), .Z(n1278) );
  XOR U1210 ( .A(n1162), .B(n1281), .Z(n1155) );
  IV U1211 ( .A(n1161), .Z(n1281) );
  XNOR U1212 ( .A(n1158), .B(n1282), .Z(n1161) );
  XOR U1213 ( .A(n1283), .B(n1284), .Z(n1158) );
  ANDN U1214 ( .A(n1285), .B(n1286), .Z(n1284) );
  XNOR U1215 ( .A(n1283), .B(n1287), .Z(n1285) );
  XOR U1216 ( .A(n1169), .B(n1288), .Z(n1162) );
  IV U1217 ( .A(n1168), .Z(n1288) );
  XNOR U1218 ( .A(n1165), .B(n1289), .Z(n1168) );
  XOR U1219 ( .A(n1290), .B(n1291), .Z(n1165) );
  ANDN U1220 ( .A(n1292), .B(n1293), .Z(n1291) );
  XNOR U1221 ( .A(n1290), .B(n1294), .Z(n1292) );
  XOR U1222 ( .A(n1176), .B(n1295), .Z(n1169) );
  IV U1223 ( .A(n1175), .Z(n1295) );
  XNOR U1224 ( .A(n1172), .B(n1296), .Z(n1175) );
  XOR U1225 ( .A(n1297), .B(n1298), .Z(n1172) );
  ANDN U1226 ( .A(n1299), .B(n1300), .Z(n1298) );
  XNOR U1227 ( .A(n1297), .B(n1301), .Z(n1299) );
  XOR U1228 ( .A(n1183), .B(n1302), .Z(n1176) );
  IV U1229 ( .A(n1182), .Z(n1302) );
  XNOR U1230 ( .A(n1179), .B(n1303), .Z(n1182) );
  XOR U1231 ( .A(n1304), .B(n1305), .Z(n1179) );
  ANDN U1232 ( .A(n1306), .B(n1307), .Z(n1305) );
  XNOR U1233 ( .A(n1304), .B(n1308), .Z(n1306) );
  XOR U1234 ( .A(n1190), .B(n1309), .Z(n1183) );
  IV U1235 ( .A(n1189), .Z(n1309) );
  XNOR U1236 ( .A(n1186), .B(n1310), .Z(n1189) );
  XOR U1237 ( .A(n1311), .B(n1312), .Z(n1186) );
  ANDN U1238 ( .A(n1313), .B(n1314), .Z(n1312) );
  XNOR U1239 ( .A(n1311), .B(n1315), .Z(n1313) );
  XOR U1240 ( .A(n1196), .B(n1316), .Z(n1190) );
  IV U1241 ( .A(n1195), .Z(n1316) );
  XNOR U1242 ( .A(n1192), .B(n1310), .Z(n1195) );
  AND U1243 ( .A(n1448), .B(n1185), .Z(n1310) );
  XOR U1244 ( .A(n1317), .B(n1318), .Z(n1192) );
  ANDN U1245 ( .A(n1319), .B(n1320), .Z(n1318) );
  XNOR U1246 ( .A(n1317), .B(n1321), .Z(n1319) );
  XOR U1247 ( .A(n1202), .B(n1322), .Z(n1196) );
  IV U1248 ( .A(n1201), .Z(n1322) );
  XNOR U1249 ( .A(n1198), .B(n1303), .Z(n1201) );
  AND U1250 ( .A(n1737), .B(n948), .Z(n1303) );
  XOR U1251 ( .A(n1323), .B(n1324), .Z(n1198) );
  ANDN U1252 ( .A(n1325), .B(n1326), .Z(n1324) );
  XNOR U1253 ( .A(n1323), .B(n1327), .Z(n1325) );
  XOR U1254 ( .A(n1208), .B(n1328), .Z(n1202) );
  IV U1255 ( .A(n1207), .Z(n1328) );
  XNOR U1256 ( .A(n1204), .B(n1296), .Z(n1207) );
  AND U1257 ( .A(n2053), .B(n736), .Z(n1296) );
  XOR U1258 ( .A(n1329), .B(n1330), .Z(n1204) );
  ANDN U1259 ( .A(n1331), .B(n1332), .Z(n1330) );
  XNOR U1260 ( .A(n1329), .B(n1333), .Z(n1331) );
  XOR U1261 ( .A(n1214), .B(n1334), .Z(n1208) );
  IV U1262 ( .A(n1213), .Z(n1334) );
  XNOR U1263 ( .A(n1210), .B(n1289), .Z(n1213) );
  AND U1264 ( .A(n2396), .B(n552), .Z(n1289) );
  XOR U1265 ( .A(n1335), .B(n1336), .Z(n1210) );
  ANDN U1266 ( .A(n1337), .B(n1338), .Z(n1336) );
  XNOR U1267 ( .A(n1335), .B(n1339), .Z(n1337) );
  XOR U1268 ( .A(n1220), .B(n1340), .Z(n1214) );
  IV U1269 ( .A(n1219), .Z(n1340) );
  XNOR U1270 ( .A(n1216), .B(n1282), .Z(n1219) );
  AND U1271 ( .A(n2765), .B(n395), .Z(n1282) );
  XOR U1272 ( .A(n1341), .B(n1342), .Z(n1216) );
  ANDN U1273 ( .A(n1343), .B(n1344), .Z(n1342) );
  XNOR U1274 ( .A(n1341), .B(n1345), .Z(n1343) );
  XOR U1275 ( .A(n1226), .B(n1346), .Z(n1220) );
  IV U1276 ( .A(n1225), .Z(n1346) );
  XNOR U1277 ( .A(n1222), .B(n1275), .Z(n1225) );
  AND U1278 ( .A(n3166), .B(n264), .Z(n1275) );
  XOR U1279 ( .A(n1347), .B(n1348), .Z(n1222) );
  ANDN U1280 ( .A(n1349), .B(n1350), .Z(n1348) );
  XNOR U1281 ( .A(n1347), .B(n1351), .Z(n1349) );
  XOR U1282 ( .A(n1232), .B(n1352), .Z(n1226) );
  IV U1283 ( .A(n1231), .Z(n1352) );
  XNOR U1284 ( .A(n1228), .B(n1268), .Z(n1231) );
  AND U1285 ( .A(n3593), .B(n159), .Z(n1268) );
  XOR U1286 ( .A(n1353), .B(n1354), .Z(n1228) );
  ANDN U1287 ( .A(n1355), .B(n1356), .Z(n1354) );
  XNOR U1288 ( .A(n1353), .B(n1357), .Z(n1355) );
  XOR U1289 ( .A(n1239), .B(n1358), .Z(n1232) );
  IV U1290 ( .A(n1238), .Z(n1358) );
  XNOR U1291 ( .A(n1235), .B(n1261), .Z(n1238) );
  AND U1292 ( .A(n4046), .B(n80), .Z(n1261) );
  XOR U1293 ( .A(n1359), .B(n1360), .Z(n1235) );
  ANDN U1294 ( .A(n1361), .B(n1362), .Z(n1360) );
  XNOR U1295 ( .A(n1359), .B(n1363), .Z(n1361) );
  XOR U1296 ( .A(n1244), .B(n1364), .Z(n1239) );
  IV U1297 ( .A(n1243), .Z(n1364) );
  XNOR U1298 ( .A(n1240), .B(n1365), .Z(n1243) );
  AND U1299 ( .A(n42), .B(n4525), .Z(n1365) );
  XOR U1300 ( .A(n1366), .B(n1367), .Z(n1240) );
  ANDN U1301 ( .A(n1368), .B(n1369), .Z(n1367) );
  XNOR U1302 ( .A(n1366), .B(n1370), .Z(n1368) );
  XNOR U1303 ( .A(n1371), .B(n1372), .Z(n1244) );
  ANDN U1304 ( .A(n1373), .B(n1374), .Z(n1372) );
  XNOR U1305 ( .A(n1371), .B(n1375), .Z(n1373) );
  XNOR U1306 ( .A(n1252), .B(n1245), .Z(n1259) );
  XOR U1307 ( .A(n1376), .B(n1377), .Z(n1245) );
  AND U1308 ( .A(n1378), .B(n1379), .Z(n1377) );
  XNOR U1309 ( .A(n9), .B(n1376), .Z(n1379) );
  XOR U1310 ( .A(n1250), .B(n1380), .Z(n1252) );
  ANDN U1311 ( .A(n4525), .B(n43), .Z(n1380) );
  XOR U1312 ( .A(n1381), .B(n1382), .Z(n1250) );
  AND U1313 ( .A(n1383), .B(n1384), .Z(n1382) );
  XNOR U1314 ( .A(n1381), .B(n1385), .Z(n1384) );
  XNOR U1315 ( .A(n794), .B(n1256), .Z(n1258) );
  AND U1316 ( .A(n1386), .B(n1387), .Z(n1256) );
  NAND U1317 ( .A(n1388), .B(n1387), .Z(n1386) );
  XOR U1318 ( .A(n1389), .B(n1378), .Z(n1388) );
  XOR U1319 ( .A(n1390), .B(n1385), .Z(n1378) );
  XOR U1320 ( .A(n1266), .B(n1391), .Z(n1385) );
  IV U1321 ( .A(n1265), .Z(n1391) );
  XNOR U1322 ( .A(n1262), .B(n1392), .Z(n1265) );
  XOR U1323 ( .A(n1393), .B(n1394), .Z(n1262) );
  ANDN U1324 ( .A(n1395), .B(n1396), .Z(n1394) );
  XNOR U1325 ( .A(n1393), .B(n1397), .Z(n1395) );
  XOR U1326 ( .A(n1273), .B(n1398), .Z(n1266) );
  IV U1327 ( .A(n1272), .Z(n1398) );
  XNOR U1328 ( .A(n1269), .B(n1399), .Z(n1272) );
  XOR U1329 ( .A(n1400), .B(n1401), .Z(n1269) );
  ANDN U1330 ( .A(n1402), .B(n1403), .Z(n1401) );
  XNOR U1331 ( .A(n1400), .B(n1404), .Z(n1402) );
  XOR U1332 ( .A(n1280), .B(n1405), .Z(n1273) );
  IV U1333 ( .A(n1279), .Z(n1405) );
  XNOR U1334 ( .A(n1276), .B(n1406), .Z(n1279) );
  XOR U1335 ( .A(n1407), .B(n1408), .Z(n1276) );
  ANDN U1336 ( .A(n1409), .B(n1410), .Z(n1408) );
  XNOR U1337 ( .A(n1407), .B(n1411), .Z(n1409) );
  XOR U1338 ( .A(n1287), .B(n1412), .Z(n1280) );
  IV U1339 ( .A(n1286), .Z(n1412) );
  XNOR U1340 ( .A(n1283), .B(n1413), .Z(n1286) );
  XOR U1341 ( .A(n1414), .B(n1415), .Z(n1283) );
  ANDN U1342 ( .A(n1416), .B(n1417), .Z(n1415) );
  XNOR U1343 ( .A(n1414), .B(n1418), .Z(n1416) );
  XOR U1344 ( .A(n1294), .B(n1419), .Z(n1287) );
  IV U1345 ( .A(n1293), .Z(n1419) );
  XNOR U1346 ( .A(n1290), .B(n1420), .Z(n1293) );
  XOR U1347 ( .A(n1421), .B(n1422), .Z(n1290) );
  ANDN U1348 ( .A(n1423), .B(n1424), .Z(n1422) );
  XNOR U1349 ( .A(n1421), .B(n1425), .Z(n1423) );
  XOR U1350 ( .A(n1301), .B(n1426), .Z(n1294) );
  IV U1351 ( .A(n1300), .Z(n1426) );
  XNOR U1352 ( .A(n1297), .B(n1427), .Z(n1300) );
  XOR U1353 ( .A(n1428), .B(n1429), .Z(n1297) );
  ANDN U1354 ( .A(n1430), .B(n1431), .Z(n1429) );
  XNOR U1355 ( .A(n1428), .B(n1432), .Z(n1430) );
  XOR U1356 ( .A(n1308), .B(n1433), .Z(n1301) );
  IV U1357 ( .A(n1307), .Z(n1433) );
  XNOR U1358 ( .A(n1304), .B(n1434), .Z(n1307) );
  XOR U1359 ( .A(n1435), .B(n1436), .Z(n1304) );
  ANDN U1360 ( .A(n1437), .B(n1438), .Z(n1436) );
  XNOR U1361 ( .A(n1435), .B(n1439), .Z(n1437) );
  XOR U1362 ( .A(n1315), .B(n1440), .Z(n1308) );
  IV U1363 ( .A(n1314), .Z(n1440) );
  XNOR U1364 ( .A(n1311), .B(n1441), .Z(n1314) );
  XOR U1365 ( .A(n1442), .B(n1443), .Z(n1311) );
  ANDN U1366 ( .A(n1444), .B(n1445), .Z(n1443) );
  XNOR U1367 ( .A(n1442), .B(n1446), .Z(n1444) );
  XOR U1368 ( .A(n1321), .B(n1447), .Z(n1315) );
  IV U1369 ( .A(n1320), .Z(n1447) );
  XNOR U1370 ( .A(n1317), .B(n1448), .Z(n1320) );
  XOR U1371 ( .A(n1449), .B(n1450), .Z(n1317) );
  ANDN U1372 ( .A(n1451), .B(n1452), .Z(n1450) );
  XNOR U1373 ( .A(n1449), .B(n1453), .Z(n1451) );
  XOR U1374 ( .A(n1327), .B(n1454), .Z(n1321) );
  IV U1375 ( .A(n1326), .Z(n1454) );
  XNOR U1376 ( .A(n1323), .B(n1441), .Z(n1326) );
  AND U1377 ( .A(n1737), .B(n1185), .Z(n1441) );
  XOR U1378 ( .A(n1455), .B(n1456), .Z(n1323) );
  ANDN U1379 ( .A(n1457), .B(n1458), .Z(n1456) );
  XNOR U1380 ( .A(n1455), .B(n1459), .Z(n1457) );
  XOR U1381 ( .A(n1333), .B(n1460), .Z(n1327) );
  IV U1382 ( .A(n1332), .Z(n1460) );
  XNOR U1383 ( .A(n1329), .B(n1434), .Z(n1332) );
  AND U1384 ( .A(n2053), .B(n948), .Z(n1434) );
  XOR U1385 ( .A(n1461), .B(n1462), .Z(n1329) );
  ANDN U1386 ( .A(n1463), .B(n1464), .Z(n1462) );
  XNOR U1387 ( .A(n1461), .B(n1465), .Z(n1463) );
  XOR U1388 ( .A(n1339), .B(n1466), .Z(n1333) );
  IV U1389 ( .A(n1338), .Z(n1466) );
  XNOR U1390 ( .A(n1335), .B(n1427), .Z(n1338) );
  AND U1391 ( .A(n2396), .B(n736), .Z(n1427) );
  XOR U1392 ( .A(n1467), .B(n1468), .Z(n1335) );
  ANDN U1393 ( .A(n1469), .B(n1470), .Z(n1468) );
  XNOR U1394 ( .A(n1467), .B(n1471), .Z(n1469) );
  XOR U1395 ( .A(n1345), .B(n1472), .Z(n1339) );
  IV U1396 ( .A(n1344), .Z(n1472) );
  XNOR U1397 ( .A(n1341), .B(n1420), .Z(n1344) );
  AND U1398 ( .A(n2765), .B(n552), .Z(n1420) );
  XOR U1399 ( .A(n1473), .B(n1474), .Z(n1341) );
  ANDN U1400 ( .A(n1475), .B(n1476), .Z(n1474) );
  XNOR U1401 ( .A(n1473), .B(n1477), .Z(n1475) );
  XOR U1402 ( .A(n1351), .B(n1478), .Z(n1345) );
  IV U1403 ( .A(n1350), .Z(n1478) );
  XNOR U1404 ( .A(n1347), .B(n1413), .Z(n1350) );
  AND U1405 ( .A(n3166), .B(n395), .Z(n1413) );
  XOR U1406 ( .A(n1479), .B(n1480), .Z(n1347) );
  ANDN U1407 ( .A(n1481), .B(n1482), .Z(n1480) );
  XNOR U1408 ( .A(n1479), .B(n1483), .Z(n1481) );
  XOR U1409 ( .A(n1357), .B(n1484), .Z(n1351) );
  IV U1410 ( .A(n1356), .Z(n1484) );
  XNOR U1411 ( .A(n1353), .B(n1406), .Z(n1356) );
  AND U1412 ( .A(n3593), .B(n264), .Z(n1406) );
  XOR U1413 ( .A(n1485), .B(n1486), .Z(n1353) );
  ANDN U1414 ( .A(n1487), .B(n1488), .Z(n1486) );
  XNOR U1415 ( .A(n1485), .B(n1489), .Z(n1487) );
  XOR U1416 ( .A(n1363), .B(n1490), .Z(n1357) );
  IV U1417 ( .A(n1362), .Z(n1490) );
  XNOR U1418 ( .A(n1359), .B(n1399), .Z(n1362) );
  AND U1419 ( .A(n4046), .B(n159), .Z(n1399) );
  XOR U1420 ( .A(n1491), .B(n1492), .Z(n1359) );
  ANDN U1421 ( .A(n1493), .B(n1494), .Z(n1492) );
  XNOR U1422 ( .A(n1491), .B(n1495), .Z(n1493) );
  XOR U1423 ( .A(n1370), .B(n1496), .Z(n1363) );
  IV U1424 ( .A(n1369), .Z(n1496) );
  XNOR U1425 ( .A(n1366), .B(n1392), .Z(n1369) );
  AND U1426 ( .A(n4525), .B(n80), .Z(n1392) );
  XOR U1427 ( .A(n1497), .B(n1498), .Z(n1366) );
  ANDN U1428 ( .A(n1499), .B(n1500), .Z(n1498) );
  XNOR U1429 ( .A(n1497), .B(n1501), .Z(n1499) );
  XOR U1430 ( .A(n1375), .B(n1502), .Z(n1370) );
  IV U1431 ( .A(n1374), .Z(n1502) );
  XNOR U1432 ( .A(n1371), .B(n1503), .Z(n1374) );
  AND U1433 ( .A(n42), .B(n5030), .Z(n1503) );
  XOR U1434 ( .A(n1504), .B(n1505), .Z(n1371) );
  ANDN U1435 ( .A(n1506), .B(n1507), .Z(n1505) );
  XNOR U1436 ( .A(n1504), .B(n1508), .Z(n1506) );
  XNOR U1437 ( .A(n1509), .B(n1510), .Z(n1375) );
  ANDN U1438 ( .A(n1511), .B(n1512), .Z(n1510) );
  XNOR U1439 ( .A(n1509), .B(n1513), .Z(n1511) );
  XNOR U1440 ( .A(n1383), .B(n1376), .Z(n1390) );
  XOR U1441 ( .A(n1514), .B(n1515), .Z(n1376) );
  AND U1442 ( .A(n1516), .B(n1517), .Z(n1515) );
  XNOR U1443 ( .A(n9), .B(n1514), .Z(n1517) );
  XOR U1444 ( .A(n1381), .B(n1518), .Z(n1383) );
  ANDN U1445 ( .A(n5030), .B(n43), .Z(n1518) );
  XOR U1446 ( .A(n1519), .B(n1520), .Z(n1381) );
  AND U1447 ( .A(n1521), .B(n1522), .Z(n1520) );
  XNOR U1448 ( .A(n1519), .B(n1523), .Z(n1522) );
  XNOR U1449 ( .A(n794), .B(n1387), .Z(n1389) );
  AND U1450 ( .A(n1524), .B(n1525), .Z(n1387) );
  NAND U1451 ( .A(n1526), .B(n1525), .Z(n1524) );
  XOR U1452 ( .A(n1527), .B(n1516), .Z(n1526) );
  XOR U1453 ( .A(n1528), .B(n1523), .Z(n1516) );
  XOR U1454 ( .A(n1397), .B(n1529), .Z(n1523) );
  IV U1455 ( .A(n1396), .Z(n1529) );
  XNOR U1456 ( .A(n1393), .B(n1530), .Z(n1396) );
  XOR U1457 ( .A(n1531), .B(n1532), .Z(n1393) );
  ANDN U1458 ( .A(n1533), .B(n1534), .Z(n1532) );
  XNOR U1459 ( .A(n1531), .B(n1535), .Z(n1533) );
  XOR U1460 ( .A(n1404), .B(n1536), .Z(n1397) );
  IV U1461 ( .A(n1403), .Z(n1536) );
  XNOR U1462 ( .A(n1400), .B(n1537), .Z(n1403) );
  XOR U1463 ( .A(n1538), .B(n1539), .Z(n1400) );
  ANDN U1464 ( .A(n1540), .B(n1541), .Z(n1539) );
  XNOR U1465 ( .A(n1538), .B(n1542), .Z(n1540) );
  XOR U1466 ( .A(n1411), .B(n1543), .Z(n1404) );
  IV U1467 ( .A(n1410), .Z(n1543) );
  XNOR U1468 ( .A(n1407), .B(n1544), .Z(n1410) );
  XOR U1469 ( .A(n1545), .B(n1546), .Z(n1407) );
  ANDN U1470 ( .A(n1547), .B(n1548), .Z(n1546) );
  XNOR U1471 ( .A(n1545), .B(n1549), .Z(n1547) );
  XOR U1472 ( .A(n1418), .B(n1550), .Z(n1411) );
  IV U1473 ( .A(n1417), .Z(n1550) );
  XNOR U1474 ( .A(n1414), .B(n1551), .Z(n1417) );
  XOR U1475 ( .A(n1552), .B(n1553), .Z(n1414) );
  ANDN U1476 ( .A(n1554), .B(n1555), .Z(n1553) );
  XNOR U1477 ( .A(n1552), .B(n1556), .Z(n1554) );
  XOR U1478 ( .A(n1425), .B(n1557), .Z(n1418) );
  IV U1479 ( .A(n1424), .Z(n1557) );
  XNOR U1480 ( .A(n1421), .B(n1558), .Z(n1424) );
  XOR U1481 ( .A(n1559), .B(n1560), .Z(n1421) );
  ANDN U1482 ( .A(n1561), .B(n1562), .Z(n1560) );
  XNOR U1483 ( .A(n1559), .B(n1563), .Z(n1561) );
  XOR U1484 ( .A(n1432), .B(n1564), .Z(n1425) );
  IV U1485 ( .A(n1431), .Z(n1564) );
  XNOR U1486 ( .A(n1428), .B(n1565), .Z(n1431) );
  XOR U1487 ( .A(n1566), .B(n1567), .Z(n1428) );
  ANDN U1488 ( .A(n1568), .B(n1569), .Z(n1567) );
  XNOR U1489 ( .A(n1566), .B(n1570), .Z(n1568) );
  XOR U1490 ( .A(n1439), .B(n1571), .Z(n1432) );
  IV U1491 ( .A(n1438), .Z(n1571) );
  XNOR U1492 ( .A(n1435), .B(n1572), .Z(n1438) );
  XOR U1493 ( .A(n1573), .B(n1574), .Z(n1435) );
  ANDN U1494 ( .A(n1575), .B(n1576), .Z(n1574) );
  XNOR U1495 ( .A(n1573), .B(n1577), .Z(n1575) );
  XOR U1496 ( .A(n1446), .B(n1578), .Z(n1439) );
  IV U1497 ( .A(n1445), .Z(n1578) );
  XNOR U1498 ( .A(n1442), .B(n1579), .Z(n1445) );
  XOR U1499 ( .A(n1580), .B(n1581), .Z(n1442) );
  ANDN U1500 ( .A(n1582), .B(n1583), .Z(n1581) );
  XNOR U1501 ( .A(n1580), .B(n1584), .Z(n1582) );
  XOR U1502 ( .A(n1453), .B(n1585), .Z(n1446) );
  IV U1503 ( .A(n1452), .Z(n1585) );
  XNOR U1504 ( .A(n1449), .B(n1586), .Z(n1452) );
  XOR U1505 ( .A(n1587), .B(n1588), .Z(n1449) );
  ANDN U1506 ( .A(n1589), .B(n1590), .Z(n1588) );
  XNOR U1507 ( .A(n1587), .B(n1591), .Z(n1589) );
  XOR U1508 ( .A(n1459), .B(n1592), .Z(n1453) );
  IV U1509 ( .A(n1458), .Z(n1592) );
  XNOR U1510 ( .A(n1455), .B(n1586), .Z(n1458) );
  AND U1511 ( .A(n1737), .B(n1448), .Z(n1586) );
  XOR U1512 ( .A(n1593), .B(n1594), .Z(n1455) );
  ANDN U1513 ( .A(n1595), .B(n1596), .Z(n1594) );
  XNOR U1514 ( .A(n1593), .B(n1597), .Z(n1595) );
  XOR U1515 ( .A(n1465), .B(n1598), .Z(n1459) );
  IV U1516 ( .A(n1464), .Z(n1598) );
  XNOR U1517 ( .A(n1461), .B(n1579), .Z(n1464) );
  AND U1518 ( .A(n2053), .B(n1185), .Z(n1579) );
  XOR U1519 ( .A(n1599), .B(n1600), .Z(n1461) );
  ANDN U1520 ( .A(n1601), .B(n1602), .Z(n1600) );
  XNOR U1521 ( .A(n1599), .B(n1603), .Z(n1601) );
  XOR U1522 ( .A(n1471), .B(n1604), .Z(n1465) );
  IV U1523 ( .A(n1470), .Z(n1604) );
  XNOR U1524 ( .A(n1467), .B(n1572), .Z(n1470) );
  AND U1525 ( .A(n2396), .B(n948), .Z(n1572) );
  XOR U1526 ( .A(n1605), .B(n1606), .Z(n1467) );
  ANDN U1527 ( .A(n1607), .B(n1608), .Z(n1606) );
  XNOR U1528 ( .A(n1605), .B(n1609), .Z(n1607) );
  XOR U1529 ( .A(n1477), .B(n1610), .Z(n1471) );
  IV U1530 ( .A(n1476), .Z(n1610) );
  XNOR U1531 ( .A(n1473), .B(n1565), .Z(n1476) );
  AND U1532 ( .A(n2765), .B(n736), .Z(n1565) );
  XOR U1533 ( .A(n1611), .B(n1612), .Z(n1473) );
  ANDN U1534 ( .A(n1613), .B(n1614), .Z(n1612) );
  XNOR U1535 ( .A(n1611), .B(n1615), .Z(n1613) );
  XOR U1536 ( .A(n1483), .B(n1616), .Z(n1477) );
  IV U1537 ( .A(n1482), .Z(n1616) );
  XNOR U1538 ( .A(n1479), .B(n1558), .Z(n1482) );
  AND U1539 ( .A(n3166), .B(n552), .Z(n1558) );
  XOR U1540 ( .A(n1617), .B(n1618), .Z(n1479) );
  ANDN U1541 ( .A(n1619), .B(n1620), .Z(n1618) );
  XNOR U1542 ( .A(n1617), .B(n1621), .Z(n1619) );
  XOR U1543 ( .A(n1489), .B(n1622), .Z(n1483) );
  IV U1544 ( .A(n1488), .Z(n1622) );
  XNOR U1545 ( .A(n1485), .B(n1551), .Z(n1488) );
  AND U1546 ( .A(n3593), .B(n395), .Z(n1551) );
  XOR U1547 ( .A(n1623), .B(n1624), .Z(n1485) );
  ANDN U1548 ( .A(n1625), .B(n1626), .Z(n1624) );
  XNOR U1549 ( .A(n1623), .B(n1627), .Z(n1625) );
  XOR U1550 ( .A(n1495), .B(n1628), .Z(n1489) );
  IV U1551 ( .A(n1494), .Z(n1628) );
  XNOR U1552 ( .A(n1491), .B(n1544), .Z(n1494) );
  AND U1553 ( .A(n4046), .B(n264), .Z(n1544) );
  XOR U1554 ( .A(n1629), .B(n1630), .Z(n1491) );
  ANDN U1555 ( .A(n1631), .B(n1632), .Z(n1630) );
  XNOR U1556 ( .A(n1629), .B(n1633), .Z(n1631) );
  XOR U1557 ( .A(n1501), .B(n1634), .Z(n1495) );
  IV U1558 ( .A(n1500), .Z(n1634) );
  XNOR U1559 ( .A(n1497), .B(n1537), .Z(n1500) );
  AND U1560 ( .A(n4525), .B(n159), .Z(n1537) );
  XOR U1561 ( .A(n1635), .B(n1636), .Z(n1497) );
  ANDN U1562 ( .A(n1637), .B(n1638), .Z(n1636) );
  XNOR U1563 ( .A(n1635), .B(n1639), .Z(n1637) );
  XOR U1564 ( .A(n1508), .B(n1640), .Z(n1501) );
  IV U1565 ( .A(n1507), .Z(n1640) );
  XNOR U1566 ( .A(n1504), .B(n1530), .Z(n1507) );
  AND U1567 ( .A(n5030), .B(n80), .Z(n1530) );
  XOR U1568 ( .A(n1641), .B(n1642), .Z(n1504) );
  ANDN U1569 ( .A(n1643), .B(n1644), .Z(n1642) );
  XNOR U1570 ( .A(n1641), .B(n1645), .Z(n1643) );
  XOR U1571 ( .A(n1513), .B(n1646), .Z(n1508) );
  IV U1572 ( .A(n1512), .Z(n1646) );
  XNOR U1573 ( .A(n1509), .B(n1647), .Z(n1512) );
  AND U1574 ( .A(n42), .B(n5561), .Z(n1647) );
  XOR U1575 ( .A(n1648), .B(n1649), .Z(n1509) );
  ANDN U1576 ( .A(n1650), .B(n1651), .Z(n1649) );
  XNOR U1577 ( .A(n1648), .B(n1652), .Z(n1650) );
  XNOR U1578 ( .A(n1653), .B(n1654), .Z(n1513) );
  ANDN U1579 ( .A(n1655), .B(n1656), .Z(n1654) );
  XNOR U1580 ( .A(n1653), .B(n1657), .Z(n1655) );
  XNOR U1581 ( .A(n1521), .B(n1514), .Z(n1528) );
  XOR U1582 ( .A(n1658), .B(n1659), .Z(n1514) );
  AND U1583 ( .A(n1660), .B(n1661), .Z(n1659) );
  XNOR U1584 ( .A(n9), .B(n1658), .Z(n1661) );
  XOR U1585 ( .A(n1519), .B(n1662), .Z(n1521) );
  ANDN U1586 ( .A(n5561), .B(n43), .Z(n1662) );
  XOR U1587 ( .A(n1663), .B(n1664), .Z(n1519) );
  AND U1588 ( .A(n1665), .B(n1666), .Z(n1664) );
  XNOR U1589 ( .A(n1663), .B(n1667), .Z(n1666) );
  XNOR U1590 ( .A(n794), .B(n1525), .Z(n1527) );
  AND U1591 ( .A(n1668), .B(n1669), .Z(n1525) );
  NAND U1592 ( .A(n1670), .B(n1669), .Z(n1668) );
  XOR U1593 ( .A(n1671), .B(n1660), .Z(n1670) );
  XOR U1594 ( .A(n1672), .B(n1667), .Z(n1660) );
  XOR U1595 ( .A(n1535), .B(n1673), .Z(n1667) );
  IV U1596 ( .A(n1534), .Z(n1673) );
  XNOR U1597 ( .A(n1531), .B(n1674), .Z(n1534) );
  XOR U1598 ( .A(n1675), .B(n1676), .Z(n1531) );
  ANDN U1599 ( .A(n1677), .B(n1678), .Z(n1676) );
  XNOR U1600 ( .A(n1675), .B(n1679), .Z(n1677) );
  XOR U1601 ( .A(n1542), .B(n1680), .Z(n1535) );
  IV U1602 ( .A(n1541), .Z(n1680) );
  XNOR U1603 ( .A(n1538), .B(n1681), .Z(n1541) );
  XOR U1604 ( .A(n1682), .B(n1683), .Z(n1538) );
  ANDN U1605 ( .A(n1684), .B(n1685), .Z(n1683) );
  XNOR U1606 ( .A(n1682), .B(n1686), .Z(n1684) );
  XOR U1607 ( .A(n1549), .B(n1687), .Z(n1542) );
  IV U1608 ( .A(n1548), .Z(n1687) );
  XNOR U1609 ( .A(n1545), .B(n1688), .Z(n1548) );
  XOR U1610 ( .A(n1689), .B(n1690), .Z(n1545) );
  ANDN U1611 ( .A(n1691), .B(n1692), .Z(n1690) );
  XNOR U1612 ( .A(n1689), .B(n1693), .Z(n1691) );
  XOR U1613 ( .A(n1556), .B(n1694), .Z(n1549) );
  IV U1614 ( .A(n1555), .Z(n1694) );
  XNOR U1615 ( .A(n1552), .B(n1695), .Z(n1555) );
  XOR U1616 ( .A(n1696), .B(n1697), .Z(n1552) );
  ANDN U1617 ( .A(n1698), .B(n1699), .Z(n1697) );
  XNOR U1618 ( .A(n1696), .B(n1700), .Z(n1698) );
  XOR U1619 ( .A(n1563), .B(n1701), .Z(n1556) );
  IV U1620 ( .A(n1562), .Z(n1701) );
  XNOR U1621 ( .A(n1559), .B(n1702), .Z(n1562) );
  XOR U1622 ( .A(n1703), .B(n1704), .Z(n1559) );
  ANDN U1623 ( .A(n1705), .B(n1706), .Z(n1704) );
  XNOR U1624 ( .A(n1703), .B(n1707), .Z(n1705) );
  XOR U1625 ( .A(n1570), .B(n1708), .Z(n1563) );
  IV U1626 ( .A(n1569), .Z(n1708) );
  XNOR U1627 ( .A(n1566), .B(n1709), .Z(n1569) );
  XOR U1628 ( .A(n1710), .B(n1711), .Z(n1566) );
  ANDN U1629 ( .A(n1712), .B(n1713), .Z(n1711) );
  XNOR U1630 ( .A(n1710), .B(n1714), .Z(n1712) );
  XOR U1631 ( .A(n1577), .B(n1715), .Z(n1570) );
  IV U1632 ( .A(n1576), .Z(n1715) );
  XNOR U1633 ( .A(n1573), .B(n1716), .Z(n1576) );
  XOR U1634 ( .A(n1717), .B(n1718), .Z(n1573) );
  ANDN U1635 ( .A(n1719), .B(n1720), .Z(n1718) );
  XNOR U1636 ( .A(n1717), .B(n1721), .Z(n1719) );
  XOR U1637 ( .A(n1584), .B(n1722), .Z(n1577) );
  IV U1638 ( .A(n1583), .Z(n1722) );
  XNOR U1639 ( .A(n1580), .B(n1723), .Z(n1583) );
  XOR U1640 ( .A(n1724), .B(n1725), .Z(n1580) );
  ANDN U1641 ( .A(n1726), .B(n1727), .Z(n1725) );
  XNOR U1642 ( .A(n1724), .B(n1728), .Z(n1726) );
  XOR U1643 ( .A(n1591), .B(n1729), .Z(n1584) );
  IV U1644 ( .A(n1590), .Z(n1729) );
  XNOR U1645 ( .A(n1587), .B(n1730), .Z(n1590) );
  XOR U1646 ( .A(n1731), .B(n1732), .Z(n1587) );
  ANDN U1647 ( .A(n1733), .B(n1734), .Z(n1732) );
  XNOR U1648 ( .A(n1731), .B(n1735), .Z(n1733) );
  XOR U1649 ( .A(n1597), .B(n1736), .Z(n1591) );
  IV U1650 ( .A(n1596), .Z(n1736) );
  XNOR U1651 ( .A(n1593), .B(n1737), .Z(n1596) );
  XOR U1652 ( .A(n1738), .B(n1739), .Z(n1593) );
  ANDN U1653 ( .A(n1740), .B(n1741), .Z(n1739) );
  XNOR U1654 ( .A(n1738), .B(n1742), .Z(n1740) );
  XOR U1655 ( .A(n1603), .B(n1743), .Z(n1597) );
  IV U1656 ( .A(n1602), .Z(n1743) );
  XNOR U1657 ( .A(n1599), .B(n1730), .Z(n1602) );
  AND U1658 ( .A(n2053), .B(n1448), .Z(n1730) );
  XOR U1659 ( .A(n1744), .B(n1745), .Z(n1599) );
  ANDN U1660 ( .A(n1746), .B(n1747), .Z(n1745) );
  XNOR U1661 ( .A(n1744), .B(n1748), .Z(n1746) );
  XOR U1662 ( .A(n1609), .B(n1749), .Z(n1603) );
  IV U1663 ( .A(n1608), .Z(n1749) );
  XNOR U1664 ( .A(n1605), .B(n1723), .Z(n1608) );
  AND U1665 ( .A(n2396), .B(n1185), .Z(n1723) );
  XOR U1666 ( .A(n1750), .B(n1751), .Z(n1605) );
  ANDN U1667 ( .A(n1752), .B(n1753), .Z(n1751) );
  XNOR U1668 ( .A(n1750), .B(n1754), .Z(n1752) );
  XOR U1669 ( .A(n1615), .B(n1755), .Z(n1609) );
  IV U1670 ( .A(n1614), .Z(n1755) );
  XNOR U1671 ( .A(n1611), .B(n1716), .Z(n1614) );
  AND U1672 ( .A(n2765), .B(n948), .Z(n1716) );
  XOR U1673 ( .A(n1756), .B(n1757), .Z(n1611) );
  ANDN U1674 ( .A(n1758), .B(n1759), .Z(n1757) );
  XNOR U1675 ( .A(n1756), .B(n1760), .Z(n1758) );
  XOR U1676 ( .A(n1621), .B(n1761), .Z(n1615) );
  IV U1677 ( .A(n1620), .Z(n1761) );
  XNOR U1678 ( .A(n1617), .B(n1709), .Z(n1620) );
  AND U1679 ( .A(n3166), .B(n736), .Z(n1709) );
  XOR U1680 ( .A(n1762), .B(n1763), .Z(n1617) );
  ANDN U1681 ( .A(n1764), .B(n1765), .Z(n1763) );
  XNOR U1682 ( .A(n1762), .B(n1766), .Z(n1764) );
  XOR U1683 ( .A(n1627), .B(n1767), .Z(n1621) );
  IV U1684 ( .A(n1626), .Z(n1767) );
  XNOR U1685 ( .A(n1623), .B(n1702), .Z(n1626) );
  AND U1686 ( .A(n3593), .B(n552), .Z(n1702) );
  XOR U1687 ( .A(n1768), .B(n1769), .Z(n1623) );
  ANDN U1688 ( .A(n1770), .B(n1771), .Z(n1769) );
  XNOR U1689 ( .A(n1768), .B(n1772), .Z(n1770) );
  XOR U1690 ( .A(n1633), .B(n1773), .Z(n1627) );
  IV U1691 ( .A(n1632), .Z(n1773) );
  XNOR U1692 ( .A(n1629), .B(n1695), .Z(n1632) );
  AND U1693 ( .A(n4046), .B(n395), .Z(n1695) );
  XOR U1694 ( .A(n1774), .B(n1775), .Z(n1629) );
  ANDN U1695 ( .A(n1776), .B(n1777), .Z(n1775) );
  XNOR U1696 ( .A(n1774), .B(n1778), .Z(n1776) );
  XOR U1697 ( .A(n1639), .B(n1779), .Z(n1633) );
  IV U1698 ( .A(n1638), .Z(n1779) );
  XNOR U1699 ( .A(n1635), .B(n1688), .Z(n1638) );
  AND U1700 ( .A(n4525), .B(n264), .Z(n1688) );
  XOR U1701 ( .A(n1780), .B(n1781), .Z(n1635) );
  ANDN U1702 ( .A(n1782), .B(n1783), .Z(n1781) );
  XNOR U1703 ( .A(n1780), .B(n1784), .Z(n1782) );
  XOR U1704 ( .A(n1645), .B(n1785), .Z(n1639) );
  IV U1705 ( .A(n1644), .Z(n1785) );
  XNOR U1706 ( .A(n1641), .B(n1681), .Z(n1644) );
  AND U1707 ( .A(n5030), .B(n159), .Z(n1681) );
  XOR U1708 ( .A(n1786), .B(n1787), .Z(n1641) );
  ANDN U1709 ( .A(n1788), .B(n1789), .Z(n1787) );
  XNOR U1710 ( .A(n1786), .B(n1790), .Z(n1788) );
  XOR U1711 ( .A(n1652), .B(n1791), .Z(n1645) );
  IV U1712 ( .A(n1651), .Z(n1791) );
  XNOR U1713 ( .A(n1648), .B(n1674), .Z(n1651) );
  AND U1714 ( .A(n5561), .B(n80), .Z(n1674) );
  XOR U1715 ( .A(n1792), .B(n1793), .Z(n1648) );
  ANDN U1716 ( .A(n1794), .B(n1795), .Z(n1793) );
  XNOR U1717 ( .A(n1792), .B(n1796), .Z(n1794) );
  XOR U1718 ( .A(n1657), .B(n1797), .Z(n1652) );
  IV U1719 ( .A(n1656), .Z(n1797) );
  XNOR U1720 ( .A(n1653), .B(n1798), .Z(n1656) );
  AND U1721 ( .A(n42), .B(n6118), .Z(n1798) );
  XOR U1722 ( .A(n1799), .B(n1800), .Z(n1653) );
  ANDN U1723 ( .A(n1801), .B(n1802), .Z(n1800) );
  XNOR U1724 ( .A(n1799), .B(n1803), .Z(n1801) );
  XNOR U1725 ( .A(n1804), .B(n1805), .Z(n1657) );
  ANDN U1726 ( .A(n1806), .B(n1807), .Z(n1805) );
  XNOR U1727 ( .A(n1804), .B(n1808), .Z(n1806) );
  XNOR U1728 ( .A(n1665), .B(n1658), .Z(n1672) );
  XOR U1729 ( .A(n1809), .B(n1810), .Z(n1658) );
  AND U1730 ( .A(n1811), .B(n1812), .Z(n1810) );
  XNOR U1731 ( .A(n9), .B(n1809), .Z(n1812) );
  XOR U1732 ( .A(n1663), .B(n1813), .Z(n1665) );
  ANDN U1733 ( .A(n6118), .B(n43), .Z(n1813) );
  XOR U1734 ( .A(n1814), .B(n1815), .Z(n1663) );
  AND U1735 ( .A(n1816), .B(n1817), .Z(n1815) );
  XNOR U1736 ( .A(n1814), .B(n1818), .Z(n1817) );
  XNOR U1737 ( .A(n794), .B(n1669), .Z(n1671) );
  AND U1738 ( .A(n1819), .B(n1820), .Z(n1669) );
  NAND U1739 ( .A(n1821), .B(n1820), .Z(n1819) );
  XOR U1740 ( .A(n1822), .B(n1811), .Z(n1821) );
  XOR U1741 ( .A(n1823), .B(n1818), .Z(n1811) );
  XOR U1742 ( .A(n1679), .B(n1824), .Z(n1818) );
  IV U1743 ( .A(n1678), .Z(n1824) );
  XNOR U1744 ( .A(n1675), .B(n1825), .Z(n1678) );
  XOR U1745 ( .A(n1826), .B(n1827), .Z(n1675) );
  ANDN U1746 ( .A(n1828), .B(n1829), .Z(n1827) );
  XNOR U1747 ( .A(n1826), .B(n1830), .Z(n1828) );
  XOR U1748 ( .A(n1686), .B(n1831), .Z(n1679) );
  IV U1749 ( .A(n1685), .Z(n1831) );
  XNOR U1750 ( .A(n1682), .B(n1832), .Z(n1685) );
  XOR U1751 ( .A(n1833), .B(n1834), .Z(n1682) );
  ANDN U1752 ( .A(n1835), .B(n1836), .Z(n1834) );
  XNOR U1753 ( .A(n1833), .B(n1837), .Z(n1835) );
  XOR U1754 ( .A(n1693), .B(n1838), .Z(n1686) );
  IV U1755 ( .A(n1692), .Z(n1838) );
  XNOR U1756 ( .A(n1689), .B(n1839), .Z(n1692) );
  XOR U1757 ( .A(n1840), .B(n1841), .Z(n1689) );
  ANDN U1758 ( .A(n1842), .B(n1843), .Z(n1841) );
  XNOR U1759 ( .A(n1840), .B(n1844), .Z(n1842) );
  XOR U1760 ( .A(n1700), .B(n1845), .Z(n1693) );
  IV U1761 ( .A(n1699), .Z(n1845) );
  XNOR U1762 ( .A(n1696), .B(n1846), .Z(n1699) );
  XOR U1763 ( .A(n1847), .B(n1848), .Z(n1696) );
  ANDN U1764 ( .A(n1849), .B(n1850), .Z(n1848) );
  XNOR U1765 ( .A(n1847), .B(n1851), .Z(n1849) );
  XOR U1766 ( .A(n1707), .B(n1852), .Z(n1700) );
  IV U1767 ( .A(n1706), .Z(n1852) );
  XNOR U1768 ( .A(n1703), .B(n1853), .Z(n1706) );
  XOR U1769 ( .A(n1854), .B(n1855), .Z(n1703) );
  ANDN U1770 ( .A(n1856), .B(n1857), .Z(n1855) );
  XNOR U1771 ( .A(n1854), .B(n1858), .Z(n1856) );
  XOR U1772 ( .A(n1714), .B(n1859), .Z(n1707) );
  IV U1773 ( .A(n1713), .Z(n1859) );
  XNOR U1774 ( .A(n1710), .B(n1860), .Z(n1713) );
  XOR U1775 ( .A(n1861), .B(n1862), .Z(n1710) );
  ANDN U1776 ( .A(n1863), .B(n1864), .Z(n1862) );
  XNOR U1777 ( .A(n1861), .B(n1865), .Z(n1863) );
  XOR U1778 ( .A(n1721), .B(n1866), .Z(n1714) );
  IV U1779 ( .A(n1720), .Z(n1866) );
  XNOR U1780 ( .A(n1717), .B(n1867), .Z(n1720) );
  XOR U1781 ( .A(n1868), .B(n1869), .Z(n1717) );
  ANDN U1782 ( .A(n1870), .B(n1871), .Z(n1869) );
  XNOR U1783 ( .A(n1868), .B(n1872), .Z(n1870) );
  XOR U1784 ( .A(n1728), .B(n1873), .Z(n1721) );
  IV U1785 ( .A(n1727), .Z(n1873) );
  XNOR U1786 ( .A(n1724), .B(n1874), .Z(n1727) );
  XOR U1787 ( .A(n1875), .B(n1876), .Z(n1724) );
  ANDN U1788 ( .A(n1877), .B(n1878), .Z(n1876) );
  XNOR U1789 ( .A(n1875), .B(n1879), .Z(n1877) );
  XOR U1790 ( .A(n1735), .B(n1880), .Z(n1728) );
  IV U1791 ( .A(n1734), .Z(n1880) );
  XNOR U1792 ( .A(n1731), .B(n1881), .Z(n1734) );
  XOR U1793 ( .A(n1882), .B(n1883), .Z(n1731) );
  ANDN U1794 ( .A(n1884), .B(n1885), .Z(n1883) );
  XNOR U1795 ( .A(n1882), .B(n1886), .Z(n1884) );
  XOR U1796 ( .A(n1742), .B(n1887), .Z(n1735) );
  IV U1797 ( .A(n1741), .Z(n1887) );
  XNOR U1798 ( .A(n1738), .B(n1888), .Z(n1741) );
  XOR U1799 ( .A(n1889), .B(n1890), .Z(n1738) );
  ANDN U1800 ( .A(n1891), .B(n1892), .Z(n1890) );
  XNOR U1801 ( .A(n1889), .B(n1893), .Z(n1891) );
  XOR U1802 ( .A(n1748), .B(n1894), .Z(n1742) );
  IV U1803 ( .A(n1747), .Z(n1894) );
  XNOR U1804 ( .A(n1744), .B(n1888), .Z(n1747) );
  AND U1805 ( .A(n2053), .B(n1737), .Z(n1888) );
  XOR U1806 ( .A(n1895), .B(n1896), .Z(n1744) );
  ANDN U1807 ( .A(n1897), .B(n1898), .Z(n1896) );
  XNOR U1808 ( .A(n1895), .B(n1899), .Z(n1897) );
  XOR U1809 ( .A(n1754), .B(n1900), .Z(n1748) );
  IV U1810 ( .A(n1753), .Z(n1900) );
  XNOR U1811 ( .A(n1750), .B(n1881), .Z(n1753) );
  AND U1812 ( .A(n2396), .B(n1448), .Z(n1881) );
  XOR U1813 ( .A(n1901), .B(n1902), .Z(n1750) );
  ANDN U1814 ( .A(n1903), .B(n1904), .Z(n1902) );
  XNOR U1815 ( .A(n1901), .B(n1905), .Z(n1903) );
  XOR U1816 ( .A(n1760), .B(n1906), .Z(n1754) );
  IV U1817 ( .A(n1759), .Z(n1906) );
  XNOR U1818 ( .A(n1756), .B(n1874), .Z(n1759) );
  AND U1819 ( .A(n2765), .B(n1185), .Z(n1874) );
  XOR U1820 ( .A(n1907), .B(n1908), .Z(n1756) );
  ANDN U1821 ( .A(n1909), .B(n1910), .Z(n1908) );
  XNOR U1822 ( .A(n1907), .B(n1911), .Z(n1909) );
  XOR U1823 ( .A(n1766), .B(n1912), .Z(n1760) );
  IV U1824 ( .A(n1765), .Z(n1912) );
  XNOR U1825 ( .A(n1762), .B(n1867), .Z(n1765) );
  AND U1826 ( .A(n3166), .B(n948), .Z(n1867) );
  XOR U1827 ( .A(n1913), .B(n1914), .Z(n1762) );
  ANDN U1828 ( .A(n1915), .B(n1916), .Z(n1914) );
  XNOR U1829 ( .A(n1913), .B(n1917), .Z(n1915) );
  XOR U1830 ( .A(n1772), .B(n1918), .Z(n1766) );
  IV U1831 ( .A(n1771), .Z(n1918) );
  XNOR U1832 ( .A(n1768), .B(n1860), .Z(n1771) );
  AND U1833 ( .A(n3593), .B(n736), .Z(n1860) );
  XOR U1834 ( .A(n1919), .B(n1920), .Z(n1768) );
  ANDN U1835 ( .A(n1921), .B(n1922), .Z(n1920) );
  XNOR U1836 ( .A(n1919), .B(n1923), .Z(n1921) );
  XOR U1837 ( .A(n1778), .B(n1924), .Z(n1772) );
  IV U1838 ( .A(n1777), .Z(n1924) );
  XNOR U1839 ( .A(n1774), .B(n1853), .Z(n1777) );
  AND U1840 ( .A(n4046), .B(n552), .Z(n1853) );
  XOR U1841 ( .A(n1925), .B(n1926), .Z(n1774) );
  ANDN U1842 ( .A(n1927), .B(n1928), .Z(n1926) );
  XNOR U1843 ( .A(n1925), .B(n1929), .Z(n1927) );
  XOR U1844 ( .A(n1784), .B(n1930), .Z(n1778) );
  IV U1845 ( .A(n1783), .Z(n1930) );
  XNOR U1846 ( .A(n1780), .B(n1846), .Z(n1783) );
  AND U1847 ( .A(n4525), .B(n395), .Z(n1846) );
  XOR U1848 ( .A(n1931), .B(n1932), .Z(n1780) );
  ANDN U1849 ( .A(n1933), .B(n1934), .Z(n1932) );
  XNOR U1850 ( .A(n1931), .B(n1935), .Z(n1933) );
  XOR U1851 ( .A(n1790), .B(n1936), .Z(n1784) );
  IV U1852 ( .A(n1789), .Z(n1936) );
  XNOR U1853 ( .A(n1786), .B(n1839), .Z(n1789) );
  AND U1854 ( .A(n5030), .B(n264), .Z(n1839) );
  XOR U1855 ( .A(n1937), .B(n1938), .Z(n1786) );
  ANDN U1856 ( .A(n1939), .B(n1940), .Z(n1938) );
  XNOR U1857 ( .A(n1937), .B(n1941), .Z(n1939) );
  XOR U1858 ( .A(n1796), .B(n1942), .Z(n1790) );
  IV U1859 ( .A(n1795), .Z(n1942) );
  XNOR U1860 ( .A(n1792), .B(n1832), .Z(n1795) );
  AND U1861 ( .A(n5561), .B(n159), .Z(n1832) );
  XOR U1862 ( .A(n1943), .B(n1944), .Z(n1792) );
  ANDN U1863 ( .A(n1945), .B(n1946), .Z(n1944) );
  XNOR U1864 ( .A(n1943), .B(n1947), .Z(n1945) );
  XOR U1865 ( .A(n1803), .B(n1948), .Z(n1796) );
  IV U1866 ( .A(n1802), .Z(n1948) );
  XNOR U1867 ( .A(n1799), .B(n1825), .Z(n1802) );
  AND U1868 ( .A(n6118), .B(n80), .Z(n1825) );
  XOR U1869 ( .A(n1949), .B(n1950), .Z(n1799) );
  ANDN U1870 ( .A(n1951), .B(n1952), .Z(n1950) );
  XNOR U1871 ( .A(n1949), .B(n1953), .Z(n1951) );
  XOR U1872 ( .A(n1808), .B(n1954), .Z(n1803) );
  IV U1873 ( .A(n1807), .Z(n1954) );
  XNOR U1874 ( .A(n1804), .B(n1955), .Z(n1807) );
  AND U1875 ( .A(n42), .B(n6688), .Z(n1955) );
  XOR U1876 ( .A(n1956), .B(n1957), .Z(n1804) );
  ANDN U1877 ( .A(n1958), .B(n1959), .Z(n1957) );
  XNOR U1878 ( .A(n1956), .B(n1960), .Z(n1958) );
  XNOR U1879 ( .A(n1961), .B(n1962), .Z(n1808) );
  ANDN U1880 ( .A(n1963), .B(n1964), .Z(n1962) );
  XNOR U1881 ( .A(n1961), .B(n1965), .Z(n1963) );
  XNOR U1882 ( .A(n1816), .B(n1809), .Z(n1823) );
  XOR U1883 ( .A(n1966), .B(n1967), .Z(n1809) );
  AND U1884 ( .A(n1968), .B(n1969), .Z(n1967) );
  XNOR U1885 ( .A(n1970), .B(n1966), .Z(n1969) );
  XOR U1886 ( .A(n1814), .B(n1971), .Z(n1816) );
  ANDN U1887 ( .A(n6688), .B(n43), .Z(n1971) );
  XOR U1888 ( .A(n1972), .B(n1973), .Z(n1814) );
  AND U1889 ( .A(n1974), .B(n1975), .Z(n1973) );
  XNOR U1890 ( .A(n1972), .B(n1976), .Z(n1975) );
  XNOR U1891 ( .A(n794), .B(n1820), .Z(n1822) );
  AND U1892 ( .A(n1977), .B(n1978), .Z(n1820) );
  NAND U1893 ( .A(n1979), .B(n1978), .Z(n1977) );
  XOR U1894 ( .A(n1980), .B(n1968), .Z(n1979) );
  XOR U1895 ( .A(n1981), .B(n1976), .Z(n1968) );
  XOR U1896 ( .A(n1830), .B(n1982), .Z(n1976) );
  IV U1897 ( .A(n1829), .Z(n1982) );
  XNOR U1898 ( .A(n1826), .B(n1983), .Z(n1829) );
  XOR U1899 ( .A(n1984), .B(n1985), .Z(n1826) );
  ANDN U1900 ( .A(n1986), .B(n1987), .Z(n1985) );
  XNOR U1901 ( .A(n1984), .B(n1988), .Z(n1986) );
  XOR U1902 ( .A(n1837), .B(n1989), .Z(n1830) );
  IV U1903 ( .A(n1836), .Z(n1989) );
  XNOR U1904 ( .A(n1833), .B(n1990), .Z(n1836) );
  XOR U1905 ( .A(n1991), .B(n1992), .Z(n1833) );
  ANDN U1906 ( .A(n1993), .B(n1994), .Z(n1992) );
  XNOR U1907 ( .A(n1991), .B(n1995), .Z(n1993) );
  XOR U1908 ( .A(n1844), .B(n1996), .Z(n1837) );
  IV U1909 ( .A(n1843), .Z(n1996) );
  XNOR U1910 ( .A(n1840), .B(n1997), .Z(n1843) );
  XOR U1911 ( .A(n1998), .B(n1999), .Z(n1840) );
  ANDN U1912 ( .A(n2000), .B(n2001), .Z(n1999) );
  XNOR U1913 ( .A(n1998), .B(n2002), .Z(n2000) );
  XOR U1914 ( .A(n1851), .B(n2003), .Z(n1844) );
  IV U1915 ( .A(n1850), .Z(n2003) );
  XNOR U1916 ( .A(n1847), .B(n2004), .Z(n1850) );
  XOR U1917 ( .A(n2005), .B(n2006), .Z(n1847) );
  ANDN U1918 ( .A(n2007), .B(n2008), .Z(n2006) );
  XNOR U1919 ( .A(n2005), .B(n2009), .Z(n2007) );
  XOR U1920 ( .A(n1858), .B(n2010), .Z(n1851) );
  IV U1921 ( .A(n1857), .Z(n2010) );
  XNOR U1922 ( .A(n1854), .B(n2011), .Z(n1857) );
  XOR U1923 ( .A(n2012), .B(n2013), .Z(n1854) );
  ANDN U1924 ( .A(n2014), .B(n2015), .Z(n2013) );
  XNOR U1925 ( .A(n2012), .B(n2016), .Z(n2014) );
  XOR U1926 ( .A(n1865), .B(n2017), .Z(n1858) );
  IV U1927 ( .A(n1864), .Z(n2017) );
  XNOR U1928 ( .A(n1861), .B(n2018), .Z(n1864) );
  XOR U1929 ( .A(n2019), .B(n2020), .Z(n1861) );
  ANDN U1930 ( .A(n2021), .B(n2022), .Z(n2020) );
  XNOR U1931 ( .A(n2019), .B(n2023), .Z(n2021) );
  XOR U1932 ( .A(n1872), .B(n2024), .Z(n1865) );
  IV U1933 ( .A(n1871), .Z(n2024) );
  XNOR U1934 ( .A(n1868), .B(n2025), .Z(n1871) );
  XOR U1935 ( .A(n2026), .B(n2027), .Z(n1868) );
  ANDN U1936 ( .A(n2028), .B(n2029), .Z(n2027) );
  XNOR U1937 ( .A(n2026), .B(n2030), .Z(n2028) );
  XOR U1938 ( .A(n1879), .B(n2031), .Z(n1872) );
  IV U1939 ( .A(n1878), .Z(n2031) );
  XNOR U1940 ( .A(n1875), .B(n2032), .Z(n1878) );
  XOR U1941 ( .A(n2033), .B(n2034), .Z(n1875) );
  ANDN U1942 ( .A(n2035), .B(n2036), .Z(n2034) );
  XNOR U1943 ( .A(n2033), .B(n2037), .Z(n2035) );
  XOR U1944 ( .A(n1886), .B(n2038), .Z(n1879) );
  IV U1945 ( .A(n1885), .Z(n2038) );
  XNOR U1946 ( .A(n1882), .B(n2039), .Z(n1885) );
  XOR U1947 ( .A(n2040), .B(n2041), .Z(n1882) );
  ANDN U1948 ( .A(n2042), .B(n2043), .Z(n2041) );
  XNOR U1949 ( .A(n2040), .B(n2044), .Z(n2042) );
  XOR U1950 ( .A(n1893), .B(n2045), .Z(n1886) );
  IV U1951 ( .A(n1892), .Z(n2045) );
  XNOR U1952 ( .A(n1889), .B(n2046), .Z(n1892) );
  XOR U1953 ( .A(n2047), .B(n2048), .Z(n1889) );
  ANDN U1954 ( .A(n2049), .B(n2050), .Z(n2048) );
  XNOR U1955 ( .A(n2047), .B(n2051), .Z(n2049) );
  XOR U1956 ( .A(n1899), .B(n2052), .Z(n1893) );
  IV U1957 ( .A(n1898), .Z(n2052) );
  XNOR U1958 ( .A(n1895), .B(n2053), .Z(n1898) );
  XOR U1959 ( .A(n2054), .B(n2055), .Z(n1895) );
  ANDN U1960 ( .A(n2056), .B(n2057), .Z(n2055) );
  XNOR U1961 ( .A(n2054), .B(n2058), .Z(n2056) );
  XOR U1962 ( .A(n1905), .B(n2059), .Z(n1899) );
  IV U1963 ( .A(n1904), .Z(n2059) );
  XNOR U1964 ( .A(n1901), .B(n2046), .Z(n1904) );
  AND U1965 ( .A(n2396), .B(n1737), .Z(n2046) );
  XOR U1966 ( .A(n2060), .B(n2061), .Z(n1901) );
  ANDN U1967 ( .A(n2062), .B(n2063), .Z(n2061) );
  XNOR U1968 ( .A(n2060), .B(n2064), .Z(n2062) );
  XOR U1969 ( .A(n1911), .B(n2065), .Z(n1905) );
  IV U1970 ( .A(n1910), .Z(n2065) );
  XNOR U1971 ( .A(n1907), .B(n2039), .Z(n1910) );
  AND U1972 ( .A(n2765), .B(n1448), .Z(n2039) );
  XOR U1973 ( .A(n2066), .B(n2067), .Z(n1907) );
  ANDN U1974 ( .A(n2068), .B(n2069), .Z(n2067) );
  XNOR U1975 ( .A(n2066), .B(n2070), .Z(n2068) );
  XOR U1976 ( .A(n1917), .B(n2071), .Z(n1911) );
  IV U1977 ( .A(n1916), .Z(n2071) );
  XNOR U1978 ( .A(n1913), .B(n2032), .Z(n1916) );
  AND U1979 ( .A(n3166), .B(n1185), .Z(n2032) );
  XOR U1980 ( .A(n2072), .B(n2073), .Z(n1913) );
  ANDN U1981 ( .A(n2074), .B(n2075), .Z(n2073) );
  XNOR U1982 ( .A(n2072), .B(n2076), .Z(n2074) );
  XOR U1983 ( .A(n1923), .B(n2077), .Z(n1917) );
  IV U1984 ( .A(n1922), .Z(n2077) );
  XNOR U1985 ( .A(n1919), .B(n2025), .Z(n1922) );
  AND U1986 ( .A(n3593), .B(n948), .Z(n2025) );
  XOR U1987 ( .A(n2078), .B(n2079), .Z(n1919) );
  ANDN U1988 ( .A(n2080), .B(n2081), .Z(n2079) );
  XNOR U1989 ( .A(n2078), .B(n2082), .Z(n2080) );
  XOR U1990 ( .A(n1929), .B(n2083), .Z(n1923) );
  IV U1991 ( .A(n1928), .Z(n2083) );
  XNOR U1992 ( .A(n1925), .B(n2018), .Z(n1928) );
  AND U1993 ( .A(n4046), .B(n736), .Z(n2018) );
  XOR U1994 ( .A(n2084), .B(n2085), .Z(n1925) );
  ANDN U1995 ( .A(n2086), .B(n2087), .Z(n2085) );
  XNOR U1996 ( .A(n2084), .B(n2088), .Z(n2086) );
  XOR U1997 ( .A(n1935), .B(n2089), .Z(n1929) );
  IV U1998 ( .A(n1934), .Z(n2089) );
  XNOR U1999 ( .A(n1931), .B(n2011), .Z(n1934) );
  AND U2000 ( .A(n4525), .B(n552), .Z(n2011) );
  XOR U2001 ( .A(n2090), .B(n2091), .Z(n1931) );
  ANDN U2002 ( .A(n2092), .B(n2093), .Z(n2091) );
  XNOR U2003 ( .A(n2090), .B(n2094), .Z(n2092) );
  XOR U2004 ( .A(n1941), .B(n2095), .Z(n1935) );
  IV U2005 ( .A(n1940), .Z(n2095) );
  XNOR U2006 ( .A(n1937), .B(n2004), .Z(n1940) );
  AND U2007 ( .A(n5030), .B(n395), .Z(n2004) );
  XOR U2008 ( .A(n2096), .B(n2097), .Z(n1937) );
  ANDN U2009 ( .A(n2098), .B(n2099), .Z(n2097) );
  XNOR U2010 ( .A(n2096), .B(n2100), .Z(n2098) );
  XOR U2011 ( .A(n1947), .B(n2101), .Z(n1941) );
  IV U2012 ( .A(n1946), .Z(n2101) );
  XNOR U2013 ( .A(n1943), .B(n1997), .Z(n1946) );
  AND U2014 ( .A(n5561), .B(n264), .Z(n1997) );
  XOR U2015 ( .A(n2102), .B(n2103), .Z(n1943) );
  ANDN U2016 ( .A(n2104), .B(n2105), .Z(n2103) );
  XNOR U2017 ( .A(n2102), .B(n2106), .Z(n2104) );
  XOR U2018 ( .A(n1953), .B(n2107), .Z(n1947) );
  IV U2019 ( .A(n1952), .Z(n2107) );
  XNOR U2020 ( .A(n1949), .B(n1990), .Z(n1952) );
  AND U2021 ( .A(n6118), .B(n159), .Z(n1990) );
  XOR U2022 ( .A(n2108), .B(n2109), .Z(n1949) );
  ANDN U2023 ( .A(n2110), .B(n2111), .Z(n2109) );
  XNOR U2024 ( .A(n2108), .B(n2112), .Z(n2110) );
  XOR U2025 ( .A(n1960), .B(n2113), .Z(n1953) );
  IV U2026 ( .A(n1959), .Z(n2113) );
  XNOR U2027 ( .A(n1956), .B(n1983), .Z(n1959) );
  AND U2028 ( .A(n6688), .B(n80), .Z(n1983) );
  XOR U2029 ( .A(n2114), .B(n2115), .Z(n1956) );
  ANDN U2030 ( .A(n2116), .B(n2117), .Z(n2115) );
  XNOR U2031 ( .A(n2114), .B(n2118), .Z(n2116) );
  XOR U2032 ( .A(n1965), .B(n2119), .Z(n1960) );
  IV U2033 ( .A(n1964), .Z(n2119) );
  XNOR U2034 ( .A(n1961), .B(n2120), .Z(n1964) );
  AND U2035 ( .A(n42), .B(n7241), .Z(n2120) );
  XOR U2036 ( .A(n2121), .B(n2122), .Z(n1961) );
  ANDN U2037 ( .A(n2123), .B(n2124), .Z(n2122) );
  XNOR U2038 ( .A(n2121), .B(n2125), .Z(n2123) );
  XNOR U2039 ( .A(n2126), .B(n2127), .Z(n1965) );
  ANDN U2040 ( .A(n2128), .B(n2129), .Z(n2127) );
  XNOR U2041 ( .A(n2126), .B(n2130), .Z(n2128) );
  XNOR U2042 ( .A(n1974), .B(n1966), .Z(n1981) );
  XOR U2043 ( .A(n2131), .B(n2132), .Z(n1966) );
  AND U2044 ( .A(n2133), .B(n2134), .Z(n2132) );
  XNOR U2045 ( .A(n2135), .B(n2131), .Z(n2134) );
  XOR U2046 ( .A(n1972), .B(n2136), .Z(n1974) );
  ANDN U2047 ( .A(n7241), .B(n43), .Z(n2136) );
  XOR U2048 ( .A(n2137), .B(n2138), .Z(n1972) );
  AND U2049 ( .A(n2139), .B(n2140), .Z(n2138) );
  XNOR U2050 ( .A(n2137), .B(n2141), .Z(n2140) );
  XOR U2051 ( .A(n1970), .B(n1978), .Z(n1980) );
  AND U2052 ( .A(n2142), .B(n2143), .Z(n1978) );
  NAND U2053 ( .A(n2144), .B(n2143), .Z(n2142) );
  XOR U2054 ( .A(n2145), .B(n2133), .Z(n2144) );
  XOR U2055 ( .A(n2146), .B(n2141), .Z(n2133) );
  XOR U2056 ( .A(n1988), .B(n2147), .Z(n2141) );
  IV U2057 ( .A(n1987), .Z(n2147) );
  XNOR U2058 ( .A(n1984), .B(n2148), .Z(n1987) );
  XOR U2059 ( .A(n2149), .B(n2150), .Z(n1984) );
  ANDN U2060 ( .A(n2151), .B(n2152), .Z(n2150) );
  XNOR U2061 ( .A(n2149), .B(n2153), .Z(n2151) );
  XOR U2062 ( .A(n1995), .B(n2154), .Z(n1988) );
  IV U2063 ( .A(n1994), .Z(n2154) );
  XNOR U2064 ( .A(n1991), .B(n2155), .Z(n1994) );
  XOR U2065 ( .A(n2156), .B(n2157), .Z(n1991) );
  ANDN U2066 ( .A(n2158), .B(n2159), .Z(n2157) );
  XNOR U2067 ( .A(n2156), .B(n2160), .Z(n2158) );
  XOR U2068 ( .A(n2002), .B(n2161), .Z(n1995) );
  IV U2069 ( .A(n2001), .Z(n2161) );
  XNOR U2070 ( .A(n1998), .B(n2162), .Z(n2001) );
  XOR U2071 ( .A(n2163), .B(n2164), .Z(n1998) );
  ANDN U2072 ( .A(n2165), .B(n2166), .Z(n2164) );
  XNOR U2073 ( .A(n2163), .B(n2167), .Z(n2165) );
  XOR U2074 ( .A(n2009), .B(n2168), .Z(n2002) );
  IV U2075 ( .A(n2008), .Z(n2168) );
  XNOR U2076 ( .A(n2005), .B(n2169), .Z(n2008) );
  XOR U2077 ( .A(n2170), .B(n2171), .Z(n2005) );
  ANDN U2078 ( .A(n2172), .B(n2173), .Z(n2171) );
  XNOR U2079 ( .A(n2170), .B(n2174), .Z(n2172) );
  XOR U2080 ( .A(n2016), .B(n2175), .Z(n2009) );
  IV U2081 ( .A(n2015), .Z(n2175) );
  XNOR U2082 ( .A(n2012), .B(n2176), .Z(n2015) );
  XOR U2083 ( .A(n2177), .B(n2178), .Z(n2012) );
  ANDN U2084 ( .A(n2179), .B(n2180), .Z(n2178) );
  XNOR U2085 ( .A(n2177), .B(n2181), .Z(n2179) );
  XOR U2086 ( .A(n2023), .B(n2182), .Z(n2016) );
  IV U2087 ( .A(n2022), .Z(n2182) );
  XNOR U2088 ( .A(n2019), .B(n2183), .Z(n2022) );
  XOR U2089 ( .A(n2184), .B(n2185), .Z(n2019) );
  ANDN U2090 ( .A(n2186), .B(n2187), .Z(n2185) );
  XNOR U2091 ( .A(n2184), .B(n2188), .Z(n2186) );
  XOR U2092 ( .A(n2030), .B(n2189), .Z(n2023) );
  IV U2093 ( .A(n2029), .Z(n2189) );
  XNOR U2094 ( .A(n2026), .B(n2190), .Z(n2029) );
  XOR U2095 ( .A(n2191), .B(n2192), .Z(n2026) );
  ANDN U2096 ( .A(n2193), .B(n2194), .Z(n2192) );
  XNOR U2097 ( .A(n2191), .B(n2195), .Z(n2193) );
  XOR U2098 ( .A(n2037), .B(n2196), .Z(n2030) );
  IV U2099 ( .A(n2036), .Z(n2196) );
  XNOR U2100 ( .A(n2033), .B(n2197), .Z(n2036) );
  XOR U2101 ( .A(n2198), .B(n2199), .Z(n2033) );
  ANDN U2102 ( .A(n2200), .B(n2201), .Z(n2199) );
  XNOR U2103 ( .A(n2198), .B(n2202), .Z(n2200) );
  XOR U2104 ( .A(n2044), .B(n2203), .Z(n2037) );
  IV U2105 ( .A(n2043), .Z(n2203) );
  XNOR U2106 ( .A(n2040), .B(n2204), .Z(n2043) );
  XOR U2107 ( .A(n2205), .B(n2206), .Z(n2040) );
  ANDN U2108 ( .A(n2207), .B(n2208), .Z(n2206) );
  XNOR U2109 ( .A(n2205), .B(n2209), .Z(n2207) );
  XOR U2110 ( .A(n2051), .B(n2210), .Z(n2044) );
  IV U2111 ( .A(n2050), .Z(n2210) );
  XNOR U2112 ( .A(n2047), .B(n2211), .Z(n2050) );
  XOR U2113 ( .A(n2212), .B(n2213), .Z(n2047) );
  ANDN U2114 ( .A(n2214), .B(n2215), .Z(n2213) );
  XNOR U2115 ( .A(n2212), .B(n2216), .Z(n2214) );
  XOR U2116 ( .A(n2058), .B(n2217), .Z(n2051) );
  IV U2117 ( .A(n2057), .Z(n2217) );
  XNOR U2118 ( .A(n2054), .B(n2218), .Z(n2057) );
  XOR U2119 ( .A(n2219), .B(n2220), .Z(n2054) );
  ANDN U2120 ( .A(n2221), .B(n2222), .Z(n2220) );
  XNOR U2121 ( .A(n2219), .B(n2223), .Z(n2221) );
  XOR U2122 ( .A(n2064), .B(n2224), .Z(n2058) );
  IV U2123 ( .A(n2063), .Z(n2224) );
  XNOR U2124 ( .A(n2060), .B(n2218), .Z(n2063) );
  AND U2125 ( .A(n2396), .B(n2053), .Z(n2218) );
  XOR U2126 ( .A(n2225), .B(n2226), .Z(n2060) );
  ANDN U2127 ( .A(n2227), .B(n2228), .Z(n2226) );
  XNOR U2128 ( .A(n2225), .B(n2229), .Z(n2227) );
  XOR U2129 ( .A(n2070), .B(n2230), .Z(n2064) );
  IV U2130 ( .A(n2069), .Z(n2230) );
  XNOR U2131 ( .A(n2066), .B(n2211), .Z(n2069) );
  AND U2132 ( .A(n2765), .B(n1737), .Z(n2211) );
  XOR U2133 ( .A(n2231), .B(n2232), .Z(n2066) );
  ANDN U2134 ( .A(n2233), .B(n2234), .Z(n2232) );
  XNOR U2135 ( .A(n2231), .B(n2235), .Z(n2233) );
  XOR U2136 ( .A(n2076), .B(n2236), .Z(n2070) );
  IV U2137 ( .A(n2075), .Z(n2236) );
  XNOR U2138 ( .A(n2072), .B(n2204), .Z(n2075) );
  AND U2139 ( .A(n3166), .B(n1448), .Z(n2204) );
  XOR U2140 ( .A(n2237), .B(n2238), .Z(n2072) );
  ANDN U2141 ( .A(n2239), .B(n2240), .Z(n2238) );
  XNOR U2142 ( .A(n2237), .B(n2241), .Z(n2239) );
  XOR U2143 ( .A(n2082), .B(n2242), .Z(n2076) );
  IV U2144 ( .A(n2081), .Z(n2242) );
  XNOR U2145 ( .A(n2078), .B(n2197), .Z(n2081) );
  AND U2146 ( .A(n3593), .B(n1185), .Z(n2197) );
  XOR U2147 ( .A(n2243), .B(n2244), .Z(n2078) );
  ANDN U2148 ( .A(n2245), .B(n2246), .Z(n2244) );
  XNOR U2149 ( .A(n2243), .B(n2247), .Z(n2245) );
  XOR U2150 ( .A(n2088), .B(n2248), .Z(n2082) );
  IV U2151 ( .A(n2087), .Z(n2248) );
  XNOR U2152 ( .A(n2084), .B(n2190), .Z(n2087) );
  AND U2153 ( .A(n4046), .B(n948), .Z(n2190) );
  XOR U2154 ( .A(n2249), .B(n2250), .Z(n2084) );
  ANDN U2155 ( .A(n2251), .B(n2252), .Z(n2250) );
  XNOR U2156 ( .A(n2249), .B(n2253), .Z(n2251) );
  XOR U2157 ( .A(n2094), .B(n2254), .Z(n2088) );
  IV U2158 ( .A(n2093), .Z(n2254) );
  XNOR U2159 ( .A(n2090), .B(n2183), .Z(n2093) );
  AND U2160 ( .A(n4525), .B(n736), .Z(n2183) );
  XOR U2161 ( .A(n2255), .B(n2256), .Z(n2090) );
  ANDN U2162 ( .A(n2257), .B(n2258), .Z(n2256) );
  XNOR U2163 ( .A(n2255), .B(n2259), .Z(n2257) );
  XOR U2164 ( .A(n2100), .B(n2260), .Z(n2094) );
  IV U2165 ( .A(n2099), .Z(n2260) );
  XNOR U2166 ( .A(n2096), .B(n2176), .Z(n2099) );
  AND U2167 ( .A(n5030), .B(n552), .Z(n2176) );
  XOR U2168 ( .A(n2261), .B(n2262), .Z(n2096) );
  ANDN U2169 ( .A(n2263), .B(n2264), .Z(n2262) );
  XNOR U2170 ( .A(n2261), .B(n2265), .Z(n2263) );
  XOR U2171 ( .A(n2106), .B(n2266), .Z(n2100) );
  IV U2172 ( .A(n2105), .Z(n2266) );
  XNOR U2173 ( .A(n2102), .B(n2169), .Z(n2105) );
  AND U2174 ( .A(n5561), .B(n395), .Z(n2169) );
  XOR U2175 ( .A(n2267), .B(n2268), .Z(n2102) );
  ANDN U2176 ( .A(n2269), .B(n2270), .Z(n2268) );
  XNOR U2177 ( .A(n2267), .B(n2271), .Z(n2269) );
  XOR U2178 ( .A(n2112), .B(n2272), .Z(n2106) );
  IV U2179 ( .A(n2111), .Z(n2272) );
  XNOR U2180 ( .A(n2108), .B(n2162), .Z(n2111) );
  AND U2181 ( .A(n6118), .B(n264), .Z(n2162) );
  XOR U2182 ( .A(n2273), .B(n2274), .Z(n2108) );
  ANDN U2183 ( .A(n2275), .B(n2276), .Z(n2274) );
  XNOR U2184 ( .A(n2273), .B(n2277), .Z(n2275) );
  XOR U2185 ( .A(n2118), .B(n2278), .Z(n2112) );
  IV U2186 ( .A(n2117), .Z(n2278) );
  XNOR U2187 ( .A(n2114), .B(n2155), .Z(n2117) );
  AND U2188 ( .A(n6688), .B(n159), .Z(n2155) );
  XOR U2189 ( .A(n2279), .B(n2280), .Z(n2114) );
  ANDN U2190 ( .A(n2281), .B(n2282), .Z(n2280) );
  XNOR U2191 ( .A(n2279), .B(n2283), .Z(n2281) );
  XOR U2192 ( .A(n2125), .B(n2284), .Z(n2118) );
  IV U2193 ( .A(n2124), .Z(n2284) );
  XNOR U2194 ( .A(n2121), .B(n2148), .Z(n2124) );
  AND U2195 ( .A(n7241), .B(n80), .Z(n2148) );
  XOR U2196 ( .A(n2285), .B(n2286), .Z(n2121) );
  ANDN U2197 ( .A(n2287), .B(n2288), .Z(n2286) );
  XNOR U2198 ( .A(n2285), .B(n2289), .Z(n2287) );
  XOR U2199 ( .A(n2130), .B(n2290), .Z(n2125) );
  IV U2200 ( .A(n2129), .Z(n2290) );
  XNOR U2201 ( .A(n2126), .B(n2291), .Z(n2129) );
  AND U2202 ( .A(n42), .B(n7770), .Z(n2291) );
  XOR U2203 ( .A(n2292), .B(n2293), .Z(n2126) );
  ANDN U2204 ( .A(n2294), .B(n2295), .Z(n2293) );
  XNOR U2205 ( .A(n2292), .B(n2296), .Z(n2294) );
  XNOR U2206 ( .A(n2297), .B(n2298), .Z(n2130) );
  ANDN U2207 ( .A(n2299), .B(n2300), .Z(n2298) );
  XNOR U2208 ( .A(n2297), .B(n2301), .Z(n2299) );
  XNOR U2209 ( .A(n2139), .B(n2131), .Z(n2146) );
  XOR U2210 ( .A(n2302), .B(n2303), .Z(n2131) );
  AND U2211 ( .A(n2304), .B(n2305), .Z(n2303) );
  XNOR U2212 ( .A(n2306), .B(n2302), .Z(n2305) );
  XOR U2213 ( .A(n2137), .B(n2307), .Z(n2139) );
  ANDN U2214 ( .A(n7770), .B(n43), .Z(n2307) );
  XOR U2215 ( .A(n2308), .B(n2309), .Z(n2137) );
  AND U2216 ( .A(n2310), .B(n2311), .Z(n2309) );
  XNOR U2217 ( .A(n2308), .B(n2312), .Z(n2311) );
  XOR U2218 ( .A(n2135), .B(n2143), .Z(n2145) );
  AND U2219 ( .A(n2313), .B(n2314), .Z(n2143) );
  NAND U2220 ( .A(n2315), .B(n2314), .Z(n2313) );
  XOR U2221 ( .A(n2316), .B(n2304), .Z(n2315) );
  XOR U2222 ( .A(n2317), .B(n2312), .Z(n2304) );
  XOR U2223 ( .A(n2153), .B(n2318), .Z(n2312) );
  IV U2224 ( .A(n2152), .Z(n2318) );
  XNOR U2225 ( .A(n2149), .B(n2319), .Z(n2152) );
  XOR U2226 ( .A(n2320), .B(n2321), .Z(n2149) );
  ANDN U2227 ( .A(n2322), .B(n2323), .Z(n2321) );
  XNOR U2228 ( .A(n2320), .B(n2324), .Z(n2322) );
  XOR U2229 ( .A(n2160), .B(n2325), .Z(n2153) );
  IV U2230 ( .A(n2159), .Z(n2325) );
  XNOR U2231 ( .A(n2156), .B(n2326), .Z(n2159) );
  XOR U2232 ( .A(n2327), .B(n2328), .Z(n2156) );
  ANDN U2233 ( .A(n2329), .B(n2330), .Z(n2328) );
  XNOR U2234 ( .A(n2327), .B(n2331), .Z(n2329) );
  XOR U2235 ( .A(n2167), .B(n2332), .Z(n2160) );
  IV U2236 ( .A(n2166), .Z(n2332) );
  XNOR U2237 ( .A(n2163), .B(n2333), .Z(n2166) );
  XOR U2238 ( .A(n2334), .B(n2335), .Z(n2163) );
  ANDN U2239 ( .A(n2336), .B(n2337), .Z(n2335) );
  XNOR U2240 ( .A(n2334), .B(n2338), .Z(n2336) );
  XOR U2241 ( .A(n2174), .B(n2339), .Z(n2167) );
  IV U2242 ( .A(n2173), .Z(n2339) );
  XNOR U2243 ( .A(n2170), .B(n2340), .Z(n2173) );
  XOR U2244 ( .A(n2341), .B(n2342), .Z(n2170) );
  ANDN U2245 ( .A(n2343), .B(n2344), .Z(n2342) );
  XNOR U2246 ( .A(n2341), .B(n2345), .Z(n2343) );
  XOR U2247 ( .A(n2181), .B(n2346), .Z(n2174) );
  IV U2248 ( .A(n2180), .Z(n2346) );
  XNOR U2249 ( .A(n2177), .B(n2347), .Z(n2180) );
  XOR U2250 ( .A(n2348), .B(n2349), .Z(n2177) );
  ANDN U2251 ( .A(n2350), .B(n2351), .Z(n2349) );
  XNOR U2252 ( .A(n2348), .B(n2352), .Z(n2350) );
  XOR U2253 ( .A(n2188), .B(n2353), .Z(n2181) );
  IV U2254 ( .A(n2187), .Z(n2353) );
  XNOR U2255 ( .A(n2184), .B(n2354), .Z(n2187) );
  XOR U2256 ( .A(n2355), .B(n2356), .Z(n2184) );
  ANDN U2257 ( .A(n2357), .B(n2358), .Z(n2356) );
  XNOR U2258 ( .A(n2355), .B(n2359), .Z(n2357) );
  XOR U2259 ( .A(n2195), .B(n2360), .Z(n2188) );
  IV U2260 ( .A(n2194), .Z(n2360) );
  XNOR U2261 ( .A(n2191), .B(n2361), .Z(n2194) );
  XOR U2262 ( .A(n2362), .B(n2363), .Z(n2191) );
  ANDN U2263 ( .A(n2364), .B(n2365), .Z(n2363) );
  XNOR U2264 ( .A(n2362), .B(n2366), .Z(n2364) );
  XOR U2265 ( .A(n2202), .B(n2367), .Z(n2195) );
  IV U2266 ( .A(n2201), .Z(n2367) );
  XNOR U2267 ( .A(n2198), .B(n2368), .Z(n2201) );
  XOR U2268 ( .A(n2369), .B(n2370), .Z(n2198) );
  ANDN U2269 ( .A(n2371), .B(n2372), .Z(n2370) );
  XNOR U2270 ( .A(n2369), .B(n2373), .Z(n2371) );
  XOR U2271 ( .A(n2209), .B(n2374), .Z(n2202) );
  IV U2272 ( .A(n2208), .Z(n2374) );
  XNOR U2273 ( .A(n2205), .B(n2375), .Z(n2208) );
  XOR U2274 ( .A(n2376), .B(n2377), .Z(n2205) );
  ANDN U2275 ( .A(n2378), .B(n2379), .Z(n2377) );
  XNOR U2276 ( .A(n2376), .B(n2380), .Z(n2378) );
  XOR U2277 ( .A(n2216), .B(n2381), .Z(n2209) );
  IV U2278 ( .A(n2215), .Z(n2381) );
  XNOR U2279 ( .A(n2212), .B(n2382), .Z(n2215) );
  XOR U2280 ( .A(n2383), .B(n2384), .Z(n2212) );
  ANDN U2281 ( .A(n2385), .B(n2386), .Z(n2384) );
  XNOR U2282 ( .A(n2383), .B(n2387), .Z(n2385) );
  XOR U2283 ( .A(n2223), .B(n2388), .Z(n2216) );
  IV U2284 ( .A(n2222), .Z(n2388) );
  XNOR U2285 ( .A(n2219), .B(n2389), .Z(n2222) );
  XOR U2286 ( .A(n2390), .B(n2391), .Z(n2219) );
  ANDN U2287 ( .A(n2392), .B(n2393), .Z(n2391) );
  XNOR U2288 ( .A(n2390), .B(n2394), .Z(n2392) );
  XOR U2289 ( .A(n2229), .B(n2395), .Z(n2223) );
  IV U2290 ( .A(n2228), .Z(n2395) );
  XNOR U2291 ( .A(n2225), .B(n2396), .Z(n2228) );
  XOR U2292 ( .A(n2397), .B(n2398), .Z(n2225) );
  ANDN U2293 ( .A(n2399), .B(n2400), .Z(n2398) );
  XNOR U2294 ( .A(n2397), .B(n2401), .Z(n2399) );
  XOR U2295 ( .A(n2235), .B(n2402), .Z(n2229) );
  IV U2296 ( .A(n2234), .Z(n2402) );
  XNOR U2297 ( .A(n2231), .B(n2389), .Z(n2234) );
  AND U2298 ( .A(n2765), .B(n2053), .Z(n2389) );
  XOR U2299 ( .A(n2403), .B(n2404), .Z(n2231) );
  ANDN U2300 ( .A(n2405), .B(n2406), .Z(n2404) );
  XNOR U2301 ( .A(n2403), .B(n2407), .Z(n2405) );
  XOR U2302 ( .A(n2241), .B(n2408), .Z(n2235) );
  IV U2303 ( .A(n2240), .Z(n2408) );
  XNOR U2304 ( .A(n2237), .B(n2382), .Z(n2240) );
  AND U2305 ( .A(n3166), .B(n1737), .Z(n2382) );
  XOR U2306 ( .A(n2409), .B(n2410), .Z(n2237) );
  ANDN U2307 ( .A(n2411), .B(n2412), .Z(n2410) );
  XNOR U2308 ( .A(n2409), .B(n2413), .Z(n2411) );
  XOR U2309 ( .A(n2247), .B(n2414), .Z(n2241) );
  IV U2310 ( .A(n2246), .Z(n2414) );
  XNOR U2311 ( .A(n2243), .B(n2375), .Z(n2246) );
  AND U2312 ( .A(n3593), .B(n1448), .Z(n2375) );
  XOR U2313 ( .A(n2415), .B(n2416), .Z(n2243) );
  ANDN U2314 ( .A(n2417), .B(n2418), .Z(n2416) );
  XNOR U2315 ( .A(n2415), .B(n2419), .Z(n2417) );
  XOR U2316 ( .A(n2253), .B(n2420), .Z(n2247) );
  IV U2317 ( .A(n2252), .Z(n2420) );
  XNOR U2318 ( .A(n2249), .B(n2368), .Z(n2252) );
  AND U2319 ( .A(n4046), .B(n1185), .Z(n2368) );
  XOR U2320 ( .A(n2421), .B(n2422), .Z(n2249) );
  ANDN U2321 ( .A(n2423), .B(n2424), .Z(n2422) );
  XNOR U2322 ( .A(n2421), .B(n2425), .Z(n2423) );
  XOR U2323 ( .A(n2259), .B(n2426), .Z(n2253) );
  IV U2324 ( .A(n2258), .Z(n2426) );
  XNOR U2325 ( .A(n2255), .B(n2361), .Z(n2258) );
  AND U2326 ( .A(n4525), .B(n948), .Z(n2361) );
  XOR U2327 ( .A(n2427), .B(n2428), .Z(n2255) );
  ANDN U2328 ( .A(n2429), .B(n2430), .Z(n2428) );
  XNOR U2329 ( .A(n2427), .B(n2431), .Z(n2429) );
  XOR U2330 ( .A(n2265), .B(n2432), .Z(n2259) );
  IV U2331 ( .A(n2264), .Z(n2432) );
  XNOR U2332 ( .A(n2261), .B(n2354), .Z(n2264) );
  AND U2333 ( .A(n5030), .B(n736), .Z(n2354) );
  XOR U2334 ( .A(n2433), .B(n2434), .Z(n2261) );
  ANDN U2335 ( .A(n2435), .B(n2436), .Z(n2434) );
  XNOR U2336 ( .A(n2433), .B(n2437), .Z(n2435) );
  XOR U2337 ( .A(n2271), .B(n2438), .Z(n2265) );
  IV U2338 ( .A(n2270), .Z(n2438) );
  XNOR U2339 ( .A(n2267), .B(n2347), .Z(n2270) );
  AND U2340 ( .A(n5561), .B(n552), .Z(n2347) );
  XOR U2341 ( .A(n2439), .B(n2440), .Z(n2267) );
  ANDN U2342 ( .A(n2441), .B(n2442), .Z(n2440) );
  XNOR U2343 ( .A(n2439), .B(n2443), .Z(n2441) );
  XOR U2344 ( .A(n2277), .B(n2444), .Z(n2271) );
  IV U2345 ( .A(n2276), .Z(n2444) );
  XNOR U2346 ( .A(n2273), .B(n2340), .Z(n2276) );
  AND U2347 ( .A(n6118), .B(n395), .Z(n2340) );
  XOR U2348 ( .A(n2445), .B(n2446), .Z(n2273) );
  ANDN U2349 ( .A(n2447), .B(n2448), .Z(n2446) );
  XNOR U2350 ( .A(n2445), .B(n2449), .Z(n2447) );
  XOR U2351 ( .A(n2283), .B(n2450), .Z(n2277) );
  IV U2352 ( .A(n2282), .Z(n2450) );
  XNOR U2353 ( .A(n2279), .B(n2333), .Z(n2282) );
  AND U2354 ( .A(n6688), .B(n264), .Z(n2333) );
  XOR U2355 ( .A(n2451), .B(n2452), .Z(n2279) );
  ANDN U2356 ( .A(n2453), .B(n2454), .Z(n2452) );
  XNOR U2357 ( .A(n2451), .B(n2455), .Z(n2453) );
  XOR U2358 ( .A(n2289), .B(n2456), .Z(n2283) );
  IV U2359 ( .A(n2288), .Z(n2456) );
  XNOR U2360 ( .A(n2285), .B(n2326), .Z(n2288) );
  AND U2361 ( .A(n7241), .B(n159), .Z(n2326) );
  XOR U2362 ( .A(n2457), .B(n2458), .Z(n2285) );
  ANDN U2363 ( .A(n2459), .B(n2460), .Z(n2458) );
  XNOR U2364 ( .A(n2457), .B(n2461), .Z(n2459) );
  XOR U2365 ( .A(n2296), .B(n2462), .Z(n2289) );
  IV U2366 ( .A(n2295), .Z(n2462) );
  XNOR U2367 ( .A(n2292), .B(n2319), .Z(n2295) );
  AND U2368 ( .A(n7770), .B(n80), .Z(n2319) );
  XOR U2369 ( .A(n2463), .B(n2464), .Z(n2292) );
  ANDN U2370 ( .A(n2465), .B(n2466), .Z(n2464) );
  XNOR U2371 ( .A(n2463), .B(n2467), .Z(n2465) );
  XOR U2372 ( .A(n2301), .B(n2468), .Z(n2296) );
  IV U2373 ( .A(n2300), .Z(n2468) );
  XNOR U2374 ( .A(n2297), .B(n2469), .Z(n2300) );
  AND U2375 ( .A(n42), .B(n8272), .Z(n2469) );
  XOR U2376 ( .A(n2470), .B(n2471), .Z(n2297) );
  ANDN U2377 ( .A(n2472), .B(n2473), .Z(n2471) );
  XNOR U2378 ( .A(n2470), .B(n2474), .Z(n2472) );
  XNOR U2379 ( .A(n2475), .B(n2476), .Z(n2301) );
  ANDN U2380 ( .A(n2477), .B(n2478), .Z(n2476) );
  XNOR U2381 ( .A(n2475), .B(n2479), .Z(n2477) );
  XNOR U2382 ( .A(n2310), .B(n2302), .Z(n2317) );
  XOR U2383 ( .A(n2480), .B(n2481), .Z(n2302) );
  AND U2384 ( .A(n2482), .B(n2483), .Z(n2481) );
  XNOR U2385 ( .A(n2484), .B(n2480), .Z(n2483) );
  XOR U2386 ( .A(n2308), .B(n2485), .Z(n2310) );
  ANDN U2387 ( .A(n8272), .B(n43), .Z(n2485) );
  XOR U2388 ( .A(n2486), .B(n2487), .Z(n2308) );
  AND U2389 ( .A(n2488), .B(n2489), .Z(n2487) );
  XNOR U2390 ( .A(n2486), .B(n2490), .Z(n2489) );
  XOR U2391 ( .A(n2306), .B(n2314), .Z(n2316) );
  AND U2392 ( .A(n2491), .B(n2492), .Z(n2314) );
  NAND U2393 ( .A(n2493), .B(n2492), .Z(n2491) );
  XOR U2394 ( .A(n2494), .B(n2482), .Z(n2493) );
  XOR U2395 ( .A(n2495), .B(n2490), .Z(n2482) );
  XOR U2396 ( .A(n2324), .B(n2496), .Z(n2490) );
  IV U2397 ( .A(n2323), .Z(n2496) );
  XNOR U2398 ( .A(n2320), .B(n2497), .Z(n2323) );
  XOR U2399 ( .A(n2498), .B(n2499), .Z(n2320) );
  ANDN U2400 ( .A(n2500), .B(n2501), .Z(n2499) );
  XNOR U2401 ( .A(n2498), .B(n2502), .Z(n2500) );
  XOR U2402 ( .A(n2331), .B(n2503), .Z(n2324) );
  IV U2403 ( .A(n2330), .Z(n2503) );
  XNOR U2404 ( .A(n2327), .B(n2504), .Z(n2330) );
  XOR U2405 ( .A(n2505), .B(n2506), .Z(n2327) );
  ANDN U2406 ( .A(n2507), .B(n2508), .Z(n2506) );
  XNOR U2407 ( .A(n2505), .B(n2509), .Z(n2507) );
  XOR U2408 ( .A(n2338), .B(n2510), .Z(n2331) );
  IV U2409 ( .A(n2337), .Z(n2510) );
  XNOR U2410 ( .A(n2334), .B(n2511), .Z(n2337) );
  XOR U2411 ( .A(n2512), .B(n2513), .Z(n2334) );
  ANDN U2412 ( .A(n2514), .B(n2515), .Z(n2513) );
  XNOR U2413 ( .A(n2512), .B(n2516), .Z(n2514) );
  XOR U2414 ( .A(n2345), .B(n2517), .Z(n2338) );
  IV U2415 ( .A(n2344), .Z(n2517) );
  XNOR U2416 ( .A(n2341), .B(n2518), .Z(n2344) );
  XOR U2417 ( .A(n2519), .B(n2520), .Z(n2341) );
  ANDN U2418 ( .A(n2521), .B(n2522), .Z(n2520) );
  XNOR U2419 ( .A(n2519), .B(n2523), .Z(n2521) );
  XOR U2420 ( .A(n2352), .B(n2524), .Z(n2345) );
  IV U2421 ( .A(n2351), .Z(n2524) );
  XNOR U2422 ( .A(n2348), .B(n2525), .Z(n2351) );
  XOR U2423 ( .A(n2526), .B(n2527), .Z(n2348) );
  ANDN U2424 ( .A(n2528), .B(n2529), .Z(n2527) );
  XNOR U2425 ( .A(n2526), .B(n2530), .Z(n2528) );
  XOR U2426 ( .A(n2359), .B(n2531), .Z(n2352) );
  IV U2427 ( .A(n2358), .Z(n2531) );
  XNOR U2428 ( .A(n2355), .B(n2532), .Z(n2358) );
  XOR U2429 ( .A(n2533), .B(n2534), .Z(n2355) );
  ANDN U2430 ( .A(n2535), .B(n2536), .Z(n2534) );
  XNOR U2431 ( .A(n2533), .B(n2537), .Z(n2535) );
  XOR U2432 ( .A(n2366), .B(n2538), .Z(n2359) );
  IV U2433 ( .A(n2365), .Z(n2538) );
  XNOR U2434 ( .A(n2362), .B(n2539), .Z(n2365) );
  XOR U2435 ( .A(n2540), .B(n2541), .Z(n2362) );
  ANDN U2436 ( .A(n2542), .B(n2543), .Z(n2541) );
  XNOR U2437 ( .A(n2540), .B(n2544), .Z(n2542) );
  XOR U2438 ( .A(n2373), .B(n2545), .Z(n2366) );
  IV U2439 ( .A(n2372), .Z(n2545) );
  XNOR U2440 ( .A(n2369), .B(n2546), .Z(n2372) );
  XOR U2441 ( .A(n2547), .B(n2548), .Z(n2369) );
  ANDN U2442 ( .A(n2549), .B(n2550), .Z(n2548) );
  XNOR U2443 ( .A(n2547), .B(n2551), .Z(n2549) );
  XOR U2444 ( .A(n2380), .B(n2552), .Z(n2373) );
  IV U2445 ( .A(n2379), .Z(n2552) );
  XNOR U2446 ( .A(n2376), .B(n2553), .Z(n2379) );
  XOR U2447 ( .A(n2554), .B(n2555), .Z(n2376) );
  ANDN U2448 ( .A(n2556), .B(n2557), .Z(n2555) );
  XNOR U2449 ( .A(n2554), .B(n2558), .Z(n2556) );
  XOR U2450 ( .A(n2387), .B(n2559), .Z(n2380) );
  IV U2451 ( .A(n2386), .Z(n2559) );
  XNOR U2452 ( .A(n2383), .B(n2560), .Z(n2386) );
  XOR U2453 ( .A(n2561), .B(n2562), .Z(n2383) );
  ANDN U2454 ( .A(n2563), .B(n2564), .Z(n2562) );
  XNOR U2455 ( .A(n2561), .B(n2565), .Z(n2563) );
  XOR U2456 ( .A(n2394), .B(n2566), .Z(n2387) );
  IV U2457 ( .A(n2393), .Z(n2566) );
  XNOR U2458 ( .A(n2390), .B(n2567), .Z(n2393) );
  XOR U2459 ( .A(n2568), .B(n2569), .Z(n2390) );
  ANDN U2460 ( .A(n2570), .B(n2571), .Z(n2569) );
  XNOR U2461 ( .A(n2568), .B(n2572), .Z(n2570) );
  XOR U2462 ( .A(n2401), .B(n2573), .Z(n2394) );
  IV U2463 ( .A(n2400), .Z(n2573) );
  XNOR U2464 ( .A(n2397), .B(n2574), .Z(n2400) );
  XOR U2465 ( .A(n2575), .B(n2576), .Z(n2397) );
  ANDN U2466 ( .A(n2577), .B(n2578), .Z(n2576) );
  XNOR U2467 ( .A(n2575), .B(n2579), .Z(n2577) );
  XOR U2468 ( .A(n2407), .B(n2580), .Z(n2401) );
  IV U2469 ( .A(n2406), .Z(n2580) );
  XNOR U2470 ( .A(n2403), .B(n2574), .Z(n2406) );
  AND U2471 ( .A(n2765), .B(n2396), .Z(n2574) );
  XOR U2472 ( .A(n2581), .B(n2582), .Z(n2403) );
  ANDN U2473 ( .A(n2583), .B(n2584), .Z(n2582) );
  XNOR U2474 ( .A(n2581), .B(n2585), .Z(n2583) );
  XOR U2475 ( .A(n2413), .B(n2586), .Z(n2407) );
  IV U2476 ( .A(n2412), .Z(n2586) );
  XNOR U2477 ( .A(n2409), .B(n2567), .Z(n2412) );
  AND U2478 ( .A(n3166), .B(n2053), .Z(n2567) );
  XOR U2479 ( .A(n2587), .B(n2588), .Z(n2409) );
  ANDN U2480 ( .A(n2589), .B(n2590), .Z(n2588) );
  XNOR U2481 ( .A(n2587), .B(n2591), .Z(n2589) );
  XOR U2482 ( .A(n2419), .B(n2592), .Z(n2413) );
  IV U2483 ( .A(n2418), .Z(n2592) );
  XNOR U2484 ( .A(n2415), .B(n2560), .Z(n2418) );
  AND U2485 ( .A(n3593), .B(n1737), .Z(n2560) );
  XOR U2486 ( .A(n2593), .B(n2594), .Z(n2415) );
  ANDN U2487 ( .A(n2595), .B(n2596), .Z(n2594) );
  XNOR U2488 ( .A(n2593), .B(n2597), .Z(n2595) );
  XOR U2489 ( .A(n2425), .B(n2598), .Z(n2419) );
  IV U2490 ( .A(n2424), .Z(n2598) );
  XNOR U2491 ( .A(n2421), .B(n2553), .Z(n2424) );
  AND U2492 ( .A(n4046), .B(n1448), .Z(n2553) );
  XOR U2493 ( .A(n2599), .B(n2600), .Z(n2421) );
  ANDN U2494 ( .A(n2601), .B(n2602), .Z(n2600) );
  XNOR U2495 ( .A(n2599), .B(n2603), .Z(n2601) );
  XOR U2496 ( .A(n2431), .B(n2604), .Z(n2425) );
  IV U2497 ( .A(n2430), .Z(n2604) );
  XNOR U2498 ( .A(n2427), .B(n2546), .Z(n2430) );
  AND U2499 ( .A(n4525), .B(n1185), .Z(n2546) );
  XOR U2500 ( .A(n2605), .B(n2606), .Z(n2427) );
  ANDN U2501 ( .A(n2607), .B(n2608), .Z(n2606) );
  XNOR U2502 ( .A(n2605), .B(n2609), .Z(n2607) );
  XOR U2503 ( .A(n2437), .B(n2610), .Z(n2431) );
  IV U2504 ( .A(n2436), .Z(n2610) );
  XNOR U2505 ( .A(n2433), .B(n2539), .Z(n2436) );
  AND U2506 ( .A(n5030), .B(n948), .Z(n2539) );
  XOR U2507 ( .A(n2611), .B(n2612), .Z(n2433) );
  ANDN U2508 ( .A(n2613), .B(n2614), .Z(n2612) );
  XNOR U2509 ( .A(n2611), .B(n2615), .Z(n2613) );
  XOR U2510 ( .A(n2443), .B(n2616), .Z(n2437) );
  IV U2511 ( .A(n2442), .Z(n2616) );
  XNOR U2512 ( .A(n2439), .B(n2532), .Z(n2442) );
  AND U2513 ( .A(n5561), .B(n736), .Z(n2532) );
  XOR U2514 ( .A(n2617), .B(n2618), .Z(n2439) );
  ANDN U2515 ( .A(n2619), .B(n2620), .Z(n2618) );
  XNOR U2516 ( .A(n2617), .B(n2621), .Z(n2619) );
  XOR U2517 ( .A(n2449), .B(n2622), .Z(n2443) );
  IV U2518 ( .A(n2448), .Z(n2622) );
  XNOR U2519 ( .A(n2445), .B(n2525), .Z(n2448) );
  AND U2520 ( .A(n6118), .B(n552), .Z(n2525) );
  XOR U2521 ( .A(n2623), .B(n2624), .Z(n2445) );
  ANDN U2522 ( .A(n2625), .B(n2626), .Z(n2624) );
  XNOR U2523 ( .A(n2623), .B(n2627), .Z(n2625) );
  XOR U2524 ( .A(n2455), .B(n2628), .Z(n2449) );
  IV U2525 ( .A(n2454), .Z(n2628) );
  XNOR U2526 ( .A(n2451), .B(n2518), .Z(n2454) );
  AND U2527 ( .A(n6688), .B(n395), .Z(n2518) );
  XOR U2528 ( .A(n2629), .B(n2630), .Z(n2451) );
  ANDN U2529 ( .A(n2631), .B(n2632), .Z(n2630) );
  XNOR U2530 ( .A(n2629), .B(n2633), .Z(n2631) );
  XOR U2531 ( .A(n2461), .B(n2634), .Z(n2455) );
  IV U2532 ( .A(n2460), .Z(n2634) );
  XNOR U2533 ( .A(n2457), .B(n2511), .Z(n2460) );
  AND U2534 ( .A(n7241), .B(n264), .Z(n2511) );
  XOR U2535 ( .A(n2635), .B(n2636), .Z(n2457) );
  ANDN U2536 ( .A(n2637), .B(n2638), .Z(n2636) );
  XNOR U2537 ( .A(n2635), .B(n2639), .Z(n2637) );
  XOR U2538 ( .A(n2467), .B(n2640), .Z(n2461) );
  IV U2539 ( .A(n2466), .Z(n2640) );
  XNOR U2540 ( .A(n2463), .B(n2504), .Z(n2466) );
  AND U2541 ( .A(n7770), .B(n159), .Z(n2504) );
  XOR U2542 ( .A(n2641), .B(n2642), .Z(n2463) );
  ANDN U2543 ( .A(n2643), .B(n2644), .Z(n2642) );
  XNOR U2544 ( .A(n2641), .B(n2645), .Z(n2643) );
  XOR U2545 ( .A(n2474), .B(n2646), .Z(n2467) );
  IV U2546 ( .A(n2473), .Z(n2646) );
  XNOR U2547 ( .A(n2470), .B(n2497), .Z(n2473) );
  AND U2548 ( .A(n8272), .B(n80), .Z(n2497) );
  XOR U2549 ( .A(n2647), .B(n2648), .Z(n2470) );
  ANDN U2550 ( .A(n2649), .B(n2650), .Z(n2648) );
  XNOR U2551 ( .A(n2647), .B(n2651), .Z(n2649) );
  XOR U2552 ( .A(n2479), .B(n2652), .Z(n2474) );
  IV U2553 ( .A(n2478), .Z(n2652) );
  XNOR U2554 ( .A(n2475), .B(n2653), .Z(n2478) );
  AND U2555 ( .A(n42), .B(n8748), .Z(n2653) );
  XOR U2556 ( .A(n2654), .B(n2655), .Z(n2475) );
  ANDN U2557 ( .A(n2656), .B(n2657), .Z(n2655) );
  XNOR U2558 ( .A(n2654), .B(n2658), .Z(n2656) );
  XNOR U2559 ( .A(n2659), .B(n2660), .Z(n2479) );
  ANDN U2560 ( .A(n2661), .B(n2662), .Z(n2660) );
  XNOR U2561 ( .A(n2659), .B(n2663), .Z(n2661) );
  XNOR U2562 ( .A(n2488), .B(n2480), .Z(n2495) );
  XOR U2563 ( .A(n2664), .B(n2665), .Z(n2480) );
  AND U2564 ( .A(n2666), .B(n2667), .Z(n2665) );
  XNOR U2565 ( .A(n2668), .B(n2664), .Z(n2667) );
  XOR U2566 ( .A(n2486), .B(n2669), .Z(n2488) );
  ANDN U2567 ( .A(n8748), .B(n43), .Z(n2669) );
  XOR U2568 ( .A(n2670), .B(n2671), .Z(n2486) );
  AND U2569 ( .A(n2672), .B(n2673), .Z(n2671) );
  XNOR U2570 ( .A(n2670), .B(n2674), .Z(n2673) );
  XOR U2571 ( .A(n2484), .B(n2492), .Z(n2494) );
  XOR U2572 ( .A(n2675), .B(n2676), .Z(n2492) );
  AND U2573 ( .A(n2675), .B(n2677), .Z(n2676) );
  XOR U2574 ( .A(n2678), .B(n2666), .Z(n2677) );
  XOR U2575 ( .A(n2679), .B(n2674), .Z(n2666) );
  XOR U2576 ( .A(n2502), .B(n2680), .Z(n2674) );
  IV U2577 ( .A(n2501), .Z(n2680) );
  XNOR U2578 ( .A(n2498), .B(n2681), .Z(n2501) );
  XOR U2579 ( .A(n2682), .B(n2683), .Z(n2498) );
  ANDN U2580 ( .A(n2684), .B(n2685), .Z(n2683) );
  XNOR U2581 ( .A(n2682), .B(n2686), .Z(n2684) );
  XOR U2582 ( .A(n2509), .B(n2687), .Z(n2502) );
  IV U2583 ( .A(n2508), .Z(n2687) );
  XNOR U2584 ( .A(n2505), .B(n2688), .Z(n2508) );
  XOR U2585 ( .A(n2689), .B(n2690), .Z(n2505) );
  ANDN U2586 ( .A(n2691), .B(n2692), .Z(n2690) );
  XNOR U2587 ( .A(n2689), .B(n2693), .Z(n2691) );
  XOR U2588 ( .A(n2516), .B(n2694), .Z(n2509) );
  IV U2589 ( .A(n2515), .Z(n2694) );
  XNOR U2590 ( .A(n2512), .B(n2695), .Z(n2515) );
  XOR U2591 ( .A(n2696), .B(n2697), .Z(n2512) );
  ANDN U2592 ( .A(n2698), .B(n2699), .Z(n2697) );
  XNOR U2593 ( .A(n2696), .B(n2700), .Z(n2698) );
  XOR U2594 ( .A(n2523), .B(n2701), .Z(n2516) );
  IV U2595 ( .A(n2522), .Z(n2701) );
  XNOR U2596 ( .A(n2519), .B(n2702), .Z(n2522) );
  XOR U2597 ( .A(n2703), .B(n2704), .Z(n2519) );
  ANDN U2598 ( .A(n2705), .B(n2706), .Z(n2704) );
  XNOR U2599 ( .A(n2703), .B(n2707), .Z(n2705) );
  XOR U2600 ( .A(n2530), .B(n2708), .Z(n2523) );
  IV U2601 ( .A(n2529), .Z(n2708) );
  XNOR U2602 ( .A(n2526), .B(n2709), .Z(n2529) );
  XOR U2603 ( .A(n2710), .B(n2711), .Z(n2526) );
  ANDN U2604 ( .A(n2712), .B(n2713), .Z(n2711) );
  XNOR U2605 ( .A(n2710), .B(n2714), .Z(n2712) );
  XOR U2606 ( .A(n2537), .B(n2715), .Z(n2530) );
  IV U2607 ( .A(n2536), .Z(n2715) );
  XNOR U2608 ( .A(n2533), .B(n2716), .Z(n2536) );
  XOR U2609 ( .A(n2717), .B(n2718), .Z(n2533) );
  ANDN U2610 ( .A(n2719), .B(n2720), .Z(n2718) );
  XNOR U2611 ( .A(n2717), .B(n2721), .Z(n2719) );
  XOR U2612 ( .A(n2544), .B(n2722), .Z(n2537) );
  IV U2613 ( .A(n2543), .Z(n2722) );
  XNOR U2614 ( .A(n2540), .B(n2723), .Z(n2543) );
  XOR U2615 ( .A(n2724), .B(n2725), .Z(n2540) );
  ANDN U2616 ( .A(n2726), .B(n2727), .Z(n2725) );
  XNOR U2617 ( .A(n2724), .B(n2728), .Z(n2726) );
  XOR U2618 ( .A(n2551), .B(n2729), .Z(n2544) );
  IV U2619 ( .A(n2550), .Z(n2729) );
  XNOR U2620 ( .A(n2547), .B(n2730), .Z(n2550) );
  XOR U2621 ( .A(n2731), .B(n2732), .Z(n2547) );
  ANDN U2622 ( .A(n2733), .B(n2734), .Z(n2732) );
  XNOR U2623 ( .A(n2731), .B(n2735), .Z(n2733) );
  XOR U2624 ( .A(n2558), .B(n2736), .Z(n2551) );
  IV U2625 ( .A(n2557), .Z(n2736) );
  XNOR U2626 ( .A(n2554), .B(n2737), .Z(n2557) );
  XOR U2627 ( .A(n2738), .B(n2739), .Z(n2554) );
  ANDN U2628 ( .A(n2740), .B(n2741), .Z(n2739) );
  XNOR U2629 ( .A(n2738), .B(n2742), .Z(n2740) );
  XOR U2630 ( .A(n2565), .B(n2743), .Z(n2558) );
  IV U2631 ( .A(n2564), .Z(n2743) );
  XNOR U2632 ( .A(n2561), .B(n2744), .Z(n2564) );
  XOR U2633 ( .A(n2745), .B(n2746), .Z(n2561) );
  ANDN U2634 ( .A(n2747), .B(n2748), .Z(n2746) );
  XNOR U2635 ( .A(n2745), .B(n2749), .Z(n2747) );
  XOR U2636 ( .A(n2572), .B(n2750), .Z(n2565) );
  IV U2637 ( .A(n2571), .Z(n2750) );
  XNOR U2638 ( .A(n2568), .B(n2751), .Z(n2571) );
  XOR U2639 ( .A(n2752), .B(n2753), .Z(n2568) );
  ANDN U2640 ( .A(n2754), .B(n2755), .Z(n2753) );
  XNOR U2641 ( .A(n2752), .B(n2756), .Z(n2754) );
  XOR U2642 ( .A(n2579), .B(n2757), .Z(n2572) );
  IV U2643 ( .A(n2578), .Z(n2757) );
  XNOR U2644 ( .A(n2575), .B(n2758), .Z(n2578) );
  XOR U2645 ( .A(n2759), .B(n2760), .Z(n2575) );
  ANDN U2646 ( .A(n2761), .B(n2762), .Z(n2760) );
  XNOR U2647 ( .A(n2759), .B(n2763), .Z(n2761) );
  XOR U2648 ( .A(n2585), .B(n2764), .Z(n2579) );
  IV U2649 ( .A(n2584), .Z(n2764) );
  XNOR U2650 ( .A(n2581), .B(n2765), .Z(n2584) );
  XOR U2651 ( .A(n2766), .B(n2767), .Z(n2581) );
  ANDN U2652 ( .A(n2768), .B(n2769), .Z(n2767) );
  XNOR U2653 ( .A(n2766), .B(n2770), .Z(n2768) );
  XOR U2654 ( .A(n2591), .B(n2771), .Z(n2585) );
  IV U2655 ( .A(n2590), .Z(n2771) );
  XNOR U2656 ( .A(n2587), .B(n2758), .Z(n2590) );
  AND U2657 ( .A(n3166), .B(n2396), .Z(n2758) );
  XOR U2658 ( .A(n2772), .B(n2773), .Z(n2587) );
  ANDN U2659 ( .A(n2774), .B(n2775), .Z(n2773) );
  XNOR U2660 ( .A(n2772), .B(n2776), .Z(n2774) );
  XOR U2661 ( .A(n2597), .B(n2777), .Z(n2591) );
  IV U2662 ( .A(n2596), .Z(n2777) );
  XNOR U2663 ( .A(n2593), .B(n2751), .Z(n2596) );
  AND U2664 ( .A(n3593), .B(n2053), .Z(n2751) );
  XOR U2665 ( .A(n2778), .B(n2779), .Z(n2593) );
  ANDN U2666 ( .A(n2780), .B(n2781), .Z(n2779) );
  XNOR U2667 ( .A(n2778), .B(n2782), .Z(n2780) );
  XOR U2668 ( .A(n2603), .B(n2783), .Z(n2597) );
  IV U2669 ( .A(n2602), .Z(n2783) );
  XNOR U2670 ( .A(n2599), .B(n2744), .Z(n2602) );
  AND U2671 ( .A(n4046), .B(n1737), .Z(n2744) );
  XOR U2672 ( .A(n2784), .B(n2785), .Z(n2599) );
  ANDN U2673 ( .A(n2786), .B(n2787), .Z(n2785) );
  XNOR U2674 ( .A(n2784), .B(n2788), .Z(n2786) );
  XOR U2675 ( .A(n2609), .B(n2789), .Z(n2603) );
  IV U2676 ( .A(n2608), .Z(n2789) );
  XNOR U2677 ( .A(n2605), .B(n2737), .Z(n2608) );
  AND U2678 ( .A(n4525), .B(n1448), .Z(n2737) );
  XOR U2679 ( .A(n2790), .B(n2791), .Z(n2605) );
  ANDN U2680 ( .A(n2792), .B(n2793), .Z(n2791) );
  XNOR U2681 ( .A(n2790), .B(n2794), .Z(n2792) );
  XOR U2682 ( .A(n2615), .B(n2795), .Z(n2609) );
  IV U2683 ( .A(n2614), .Z(n2795) );
  XNOR U2684 ( .A(n2611), .B(n2730), .Z(n2614) );
  AND U2685 ( .A(n5030), .B(n1185), .Z(n2730) );
  XOR U2686 ( .A(n2796), .B(n2797), .Z(n2611) );
  ANDN U2687 ( .A(n2798), .B(n2799), .Z(n2797) );
  XNOR U2688 ( .A(n2796), .B(n2800), .Z(n2798) );
  XOR U2689 ( .A(n2621), .B(n2801), .Z(n2615) );
  IV U2690 ( .A(n2620), .Z(n2801) );
  XNOR U2691 ( .A(n2617), .B(n2723), .Z(n2620) );
  AND U2692 ( .A(n5561), .B(n948), .Z(n2723) );
  XOR U2693 ( .A(n2802), .B(n2803), .Z(n2617) );
  ANDN U2694 ( .A(n2804), .B(n2805), .Z(n2803) );
  XNOR U2695 ( .A(n2802), .B(n2806), .Z(n2804) );
  XOR U2696 ( .A(n2627), .B(n2807), .Z(n2621) );
  IV U2697 ( .A(n2626), .Z(n2807) );
  XNOR U2698 ( .A(n2623), .B(n2716), .Z(n2626) );
  AND U2699 ( .A(n6118), .B(n736), .Z(n2716) );
  XOR U2700 ( .A(n2808), .B(n2809), .Z(n2623) );
  ANDN U2701 ( .A(n2810), .B(n2811), .Z(n2809) );
  XNOR U2702 ( .A(n2808), .B(n2812), .Z(n2810) );
  XOR U2703 ( .A(n2633), .B(n2813), .Z(n2627) );
  IV U2704 ( .A(n2632), .Z(n2813) );
  XNOR U2705 ( .A(n2629), .B(n2709), .Z(n2632) );
  AND U2706 ( .A(n6688), .B(n552), .Z(n2709) );
  XOR U2707 ( .A(n2814), .B(n2815), .Z(n2629) );
  ANDN U2708 ( .A(n2816), .B(n2817), .Z(n2815) );
  XNOR U2709 ( .A(n2814), .B(n2818), .Z(n2816) );
  XOR U2710 ( .A(n2639), .B(n2819), .Z(n2633) );
  IV U2711 ( .A(n2638), .Z(n2819) );
  XNOR U2712 ( .A(n2635), .B(n2702), .Z(n2638) );
  AND U2713 ( .A(n7241), .B(n395), .Z(n2702) );
  XOR U2714 ( .A(n2820), .B(n2821), .Z(n2635) );
  ANDN U2715 ( .A(n2822), .B(n2823), .Z(n2821) );
  XNOR U2716 ( .A(n2820), .B(n2824), .Z(n2822) );
  XOR U2717 ( .A(n2645), .B(n2825), .Z(n2639) );
  IV U2718 ( .A(n2644), .Z(n2825) );
  XNOR U2719 ( .A(n2641), .B(n2695), .Z(n2644) );
  AND U2720 ( .A(n7770), .B(n264), .Z(n2695) );
  XOR U2721 ( .A(n2826), .B(n2827), .Z(n2641) );
  ANDN U2722 ( .A(n2828), .B(n2829), .Z(n2827) );
  XNOR U2723 ( .A(n2826), .B(n2830), .Z(n2828) );
  XOR U2724 ( .A(n2651), .B(n2831), .Z(n2645) );
  IV U2725 ( .A(n2650), .Z(n2831) );
  XNOR U2726 ( .A(n2647), .B(n2688), .Z(n2650) );
  AND U2727 ( .A(n8272), .B(n159), .Z(n2688) );
  XOR U2728 ( .A(n2832), .B(n2833), .Z(n2647) );
  ANDN U2729 ( .A(n2834), .B(n2835), .Z(n2833) );
  XNOR U2730 ( .A(n2832), .B(n2836), .Z(n2834) );
  XOR U2731 ( .A(n2658), .B(n2837), .Z(n2651) );
  IV U2732 ( .A(n2657), .Z(n2837) );
  XNOR U2733 ( .A(n2654), .B(n2681), .Z(n2657) );
  AND U2734 ( .A(n8748), .B(n80), .Z(n2681) );
  XOR U2735 ( .A(n2838), .B(n2839), .Z(n2654) );
  ANDN U2736 ( .A(n2840), .B(n2841), .Z(n2839) );
  XNOR U2737 ( .A(n2838), .B(n2842), .Z(n2840) );
  XOR U2738 ( .A(n2663), .B(n2843), .Z(n2658) );
  IV U2739 ( .A(n2662), .Z(n2843) );
  XNOR U2740 ( .A(n2659), .B(n2844), .Z(n2662) );
  AND U2741 ( .A(n42), .B(n9198), .Z(n2844) );
  XOR U2742 ( .A(n2845), .B(n2846), .Z(n2659) );
  ANDN U2743 ( .A(n2847), .B(n2848), .Z(n2846) );
  XNOR U2744 ( .A(n2845), .B(n2849), .Z(n2847) );
  XNOR U2745 ( .A(n2850), .B(n2851), .Z(n2663) );
  ANDN U2746 ( .A(n2852), .B(n2853), .Z(n2851) );
  XNOR U2747 ( .A(n2850), .B(n2854), .Z(n2852) );
  XNOR U2748 ( .A(n2672), .B(n2664), .Z(n2679) );
  XOR U2749 ( .A(n2855), .B(n2856), .Z(n2664) );
  AND U2750 ( .A(n2857), .B(n2858), .Z(n2856) );
  XNOR U2751 ( .A(n2859), .B(n2855), .Z(n2858) );
  XOR U2752 ( .A(n2670), .B(n2860), .Z(n2672) );
  ANDN U2753 ( .A(n9198), .B(n43), .Z(n2860) );
  XOR U2754 ( .A(n2861), .B(n2862), .Z(n2670) );
  AND U2755 ( .A(n2863), .B(n2864), .Z(n2862) );
  XNOR U2756 ( .A(n2861), .B(n2865), .Z(n2864) );
  XOR U2757 ( .A(n2668), .B(n2675), .Z(n2678) );
  XOR U2758 ( .A(n2866), .B(n2867), .Z(n2668) );
  IV U2759 ( .A(n2868), .Z(n2867) );
  XOR U2760 ( .A(n2869), .B(n2870), .Z(n2675) );
  AND U2761 ( .A(n2869), .B(n2871), .Z(n2870) );
  XOR U2762 ( .A(n2872), .B(n2857), .Z(n2871) );
  XOR U2763 ( .A(n2873), .B(n2865), .Z(n2857) );
  XOR U2764 ( .A(n2686), .B(n2874), .Z(n2865) );
  IV U2765 ( .A(n2685), .Z(n2874) );
  XNOR U2766 ( .A(n2682), .B(n2875), .Z(n2685) );
  XOR U2767 ( .A(n2876), .B(n2877), .Z(n2682) );
  ANDN U2768 ( .A(n2878), .B(n2879), .Z(n2877) );
  XNOR U2769 ( .A(n2876), .B(n2880), .Z(n2878) );
  XOR U2770 ( .A(n2693), .B(n2881), .Z(n2686) );
  IV U2771 ( .A(n2692), .Z(n2881) );
  XNOR U2772 ( .A(n2689), .B(n2882), .Z(n2692) );
  XOR U2773 ( .A(n2883), .B(n2884), .Z(n2689) );
  ANDN U2774 ( .A(n2885), .B(n2886), .Z(n2884) );
  XNOR U2775 ( .A(n2883), .B(n2887), .Z(n2885) );
  XOR U2776 ( .A(n2700), .B(n2888), .Z(n2693) );
  IV U2777 ( .A(n2699), .Z(n2888) );
  XNOR U2778 ( .A(n2696), .B(n2889), .Z(n2699) );
  XOR U2779 ( .A(n2890), .B(n2891), .Z(n2696) );
  ANDN U2780 ( .A(n2892), .B(n2893), .Z(n2891) );
  XNOR U2781 ( .A(n2890), .B(n2894), .Z(n2892) );
  XOR U2782 ( .A(n2707), .B(n2895), .Z(n2700) );
  IV U2783 ( .A(n2706), .Z(n2895) );
  XNOR U2784 ( .A(n2703), .B(n2896), .Z(n2706) );
  XOR U2785 ( .A(n2897), .B(n2898), .Z(n2703) );
  ANDN U2786 ( .A(n2899), .B(n2900), .Z(n2898) );
  XNOR U2787 ( .A(n2897), .B(n2901), .Z(n2899) );
  XOR U2788 ( .A(n2714), .B(n2902), .Z(n2707) );
  IV U2789 ( .A(n2713), .Z(n2902) );
  XNOR U2790 ( .A(n2710), .B(n2903), .Z(n2713) );
  XOR U2791 ( .A(n2904), .B(n2905), .Z(n2710) );
  ANDN U2792 ( .A(n2906), .B(n2907), .Z(n2905) );
  XNOR U2793 ( .A(n2904), .B(n2908), .Z(n2906) );
  XOR U2794 ( .A(n2721), .B(n2909), .Z(n2714) );
  IV U2795 ( .A(n2720), .Z(n2909) );
  XNOR U2796 ( .A(n2717), .B(n2910), .Z(n2720) );
  XOR U2797 ( .A(n2911), .B(n2912), .Z(n2717) );
  ANDN U2798 ( .A(n2913), .B(n2914), .Z(n2912) );
  XNOR U2799 ( .A(n2911), .B(n2915), .Z(n2913) );
  XOR U2800 ( .A(n2728), .B(n2916), .Z(n2721) );
  IV U2801 ( .A(n2727), .Z(n2916) );
  XNOR U2802 ( .A(n2724), .B(n2917), .Z(n2727) );
  XOR U2803 ( .A(n2918), .B(n2919), .Z(n2724) );
  ANDN U2804 ( .A(n2920), .B(n2921), .Z(n2919) );
  XNOR U2805 ( .A(n2918), .B(n2922), .Z(n2920) );
  XOR U2806 ( .A(n2735), .B(n2923), .Z(n2728) );
  IV U2807 ( .A(n2734), .Z(n2923) );
  XNOR U2808 ( .A(n2731), .B(n2924), .Z(n2734) );
  XOR U2809 ( .A(n2925), .B(n2926), .Z(n2731) );
  ANDN U2810 ( .A(n2927), .B(n2928), .Z(n2926) );
  XNOR U2811 ( .A(n2925), .B(n2929), .Z(n2927) );
  XOR U2812 ( .A(n2742), .B(n2930), .Z(n2735) );
  IV U2813 ( .A(n2741), .Z(n2930) );
  XNOR U2814 ( .A(n2738), .B(n2931), .Z(n2741) );
  XOR U2815 ( .A(n2932), .B(n2933), .Z(n2738) );
  ANDN U2816 ( .A(n2934), .B(n2935), .Z(n2933) );
  XNOR U2817 ( .A(n2932), .B(n2936), .Z(n2934) );
  XOR U2818 ( .A(n2749), .B(n2937), .Z(n2742) );
  IV U2819 ( .A(n2748), .Z(n2937) );
  XNOR U2820 ( .A(n2745), .B(n2938), .Z(n2748) );
  XOR U2821 ( .A(n2939), .B(n2940), .Z(n2745) );
  ANDN U2822 ( .A(n2941), .B(n2942), .Z(n2940) );
  XNOR U2823 ( .A(n2939), .B(n2943), .Z(n2941) );
  XOR U2824 ( .A(n2756), .B(n2944), .Z(n2749) );
  IV U2825 ( .A(n2755), .Z(n2944) );
  XNOR U2826 ( .A(n2752), .B(n2945), .Z(n2755) );
  XOR U2827 ( .A(n2946), .B(n2947), .Z(n2752) );
  ANDN U2828 ( .A(n2948), .B(n2949), .Z(n2947) );
  XNOR U2829 ( .A(n2946), .B(n2950), .Z(n2948) );
  XOR U2830 ( .A(n2763), .B(n2951), .Z(n2756) );
  IV U2831 ( .A(n2762), .Z(n2951) );
  XNOR U2832 ( .A(n2759), .B(n2952), .Z(n2762) );
  XOR U2833 ( .A(n2953), .B(n2954), .Z(n2759) );
  ANDN U2834 ( .A(n2955), .B(n2956), .Z(n2954) );
  XNOR U2835 ( .A(n2953), .B(n2957), .Z(n2955) );
  XOR U2836 ( .A(n2770), .B(n2958), .Z(n2763) );
  IV U2837 ( .A(n2769), .Z(n2958) );
  XNOR U2838 ( .A(n2766), .B(n2959), .Z(n2769) );
  XOR U2839 ( .A(n2960), .B(n2961), .Z(n2766) );
  ANDN U2840 ( .A(n2962), .B(n2963), .Z(n2961) );
  XNOR U2841 ( .A(n2960), .B(n2964), .Z(n2962) );
  XOR U2842 ( .A(n2776), .B(n2965), .Z(n2770) );
  IV U2843 ( .A(n2775), .Z(n2965) );
  XNOR U2844 ( .A(n2772), .B(n2959), .Z(n2775) );
  AND U2845 ( .A(n3166), .B(n2765), .Z(n2959) );
  XOR U2846 ( .A(n2966), .B(n2967), .Z(n2772) );
  ANDN U2847 ( .A(n2968), .B(n2969), .Z(n2967) );
  XNOR U2848 ( .A(n2966), .B(n2970), .Z(n2968) );
  XOR U2849 ( .A(n2782), .B(n2971), .Z(n2776) );
  IV U2850 ( .A(n2781), .Z(n2971) );
  XNOR U2851 ( .A(n2778), .B(n2952), .Z(n2781) );
  AND U2852 ( .A(n3593), .B(n2396), .Z(n2952) );
  XOR U2853 ( .A(n2972), .B(n2973), .Z(n2778) );
  ANDN U2854 ( .A(n2974), .B(n2975), .Z(n2973) );
  XNOR U2855 ( .A(n2972), .B(n2976), .Z(n2974) );
  XOR U2856 ( .A(n2788), .B(n2977), .Z(n2782) );
  IV U2857 ( .A(n2787), .Z(n2977) );
  XNOR U2858 ( .A(n2784), .B(n2945), .Z(n2787) );
  AND U2859 ( .A(n4046), .B(n2053), .Z(n2945) );
  XOR U2860 ( .A(n2978), .B(n2979), .Z(n2784) );
  ANDN U2861 ( .A(n2980), .B(n2981), .Z(n2979) );
  XNOR U2862 ( .A(n2978), .B(n2982), .Z(n2980) );
  XOR U2863 ( .A(n2794), .B(n2983), .Z(n2788) );
  IV U2864 ( .A(n2793), .Z(n2983) );
  XNOR U2865 ( .A(n2790), .B(n2938), .Z(n2793) );
  AND U2866 ( .A(n4525), .B(n1737), .Z(n2938) );
  XOR U2867 ( .A(n2984), .B(n2985), .Z(n2790) );
  ANDN U2868 ( .A(n2986), .B(n2987), .Z(n2985) );
  XNOR U2869 ( .A(n2984), .B(n2988), .Z(n2986) );
  XOR U2870 ( .A(n2800), .B(n2989), .Z(n2794) );
  IV U2871 ( .A(n2799), .Z(n2989) );
  XNOR U2872 ( .A(n2796), .B(n2931), .Z(n2799) );
  AND U2873 ( .A(n5030), .B(n1448), .Z(n2931) );
  XOR U2874 ( .A(n2990), .B(n2991), .Z(n2796) );
  ANDN U2875 ( .A(n2992), .B(n2993), .Z(n2991) );
  XNOR U2876 ( .A(n2990), .B(n2994), .Z(n2992) );
  XOR U2877 ( .A(n2806), .B(n2995), .Z(n2800) );
  IV U2878 ( .A(n2805), .Z(n2995) );
  XNOR U2879 ( .A(n2802), .B(n2924), .Z(n2805) );
  AND U2880 ( .A(n5561), .B(n1185), .Z(n2924) );
  XOR U2881 ( .A(n2996), .B(n2997), .Z(n2802) );
  ANDN U2882 ( .A(n2998), .B(n2999), .Z(n2997) );
  XNOR U2883 ( .A(n2996), .B(n3000), .Z(n2998) );
  XOR U2884 ( .A(n2812), .B(n3001), .Z(n2806) );
  IV U2885 ( .A(n2811), .Z(n3001) );
  XNOR U2886 ( .A(n2808), .B(n2917), .Z(n2811) );
  AND U2887 ( .A(n6118), .B(n948), .Z(n2917) );
  XOR U2888 ( .A(n3002), .B(n3003), .Z(n2808) );
  ANDN U2889 ( .A(n3004), .B(n3005), .Z(n3003) );
  XNOR U2890 ( .A(n3002), .B(n3006), .Z(n3004) );
  XOR U2891 ( .A(n2818), .B(n3007), .Z(n2812) );
  IV U2892 ( .A(n2817), .Z(n3007) );
  XNOR U2893 ( .A(n2814), .B(n2910), .Z(n2817) );
  AND U2894 ( .A(n6688), .B(n736), .Z(n2910) );
  XOR U2895 ( .A(n3008), .B(n3009), .Z(n2814) );
  ANDN U2896 ( .A(n3010), .B(n3011), .Z(n3009) );
  XNOR U2897 ( .A(n3008), .B(n3012), .Z(n3010) );
  XOR U2898 ( .A(n2824), .B(n3013), .Z(n2818) );
  IV U2899 ( .A(n2823), .Z(n3013) );
  XNOR U2900 ( .A(n2820), .B(n2903), .Z(n2823) );
  AND U2901 ( .A(n7241), .B(n552), .Z(n2903) );
  XOR U2902 ( .A(n3014), .B(n3015), .Z(n2820) );
  ANDN U2903 ( .A(n3016), .B(n3017), .Z(n3015) );
  XNOR U2904 ( .A(n3014), .B(n3018), .Z(n3016) );
  XOR U2905 ( .A(n2830), .B(n3019), .Z(n2824) );
  IV U2906 ( .A(n2829), .Z(n3019) );
  XNOR U2907 ( .A(n2826), .B(n2896), .Z(n2829) );
  AND U2908 ( .A(n7770), .B(n395), .Z(n2896) );
  XOR U2909 ( .A(n3020), .B(n3021), .Z(n2826) );
  ANDN U2910 ( .A(n3022), .B(n3023), .Z(n3021) );
  XNOR U2911 ( .A(n3020), .B(n3024), .Z(n3022) );
  XOR U2912 ( .A(n2836), .B(n3025), .Z(n2830) );
  IV U2913 ( .A(n2835), .Z(n3025) );
  XNOR U2914 ( .A(n2832), .B(n2889), .Z(n2835) );
  AND U2915 ( .A(n8272), .B(n264), .Z(n2889) );
  XOR U2916 ( .A(n3026), .B(n3027), .Z(n2832) );
  ANDN U2917 ( .A(n3028), .B(n3029), .Z(n3027) );
  XNOR U2918 ( .A(n3026), .B(n3030), .Z(n3028) );
  XOR U2919 ( .A(n2842), .B(n3031), .Z(n2836) );
  IV U2920 ( .A(n2841), .Z(n3031) );
  XNOR U2921 ( .A(n2838), .B(n2882), .Z(n2841) );
  AND U2922 ( .A(n8748), .B(n159), .Z(n2882) );
  XOR U2923 ( .A(n3032), .B(n3033), .Z(n2838) );
  ANDN U2924 ( .A(n3034), .B(n3035), .Z(n3033) );
  XNOR U2925 ( .A(n3032), .B(n3036), .Z(n3034) );
  XOR U2926 ( .A(n2849), .B(n3037), .Z(n2842) );
  IV U2927 ( .A(n2848), .Z(n3037) );
  XNOR U2928 ( .A(n2845), .B(n2875), .Z(n2848) );
  AND U2929 ( .A(n9198), .B(n80), .Z(n2875) );
  XOR U2930 ( .A(n3038), .B(n3039), .Z(n2845) );
  ANDN U2931 ( .A(n3040), .B(n3041), .Z(n3039) );
  XNOR U2932 ( .A(n3038), .B(n3042), .Z(n3040) );
  XOR U2933 ( .A(n2854), .B(n3043), .Z(n2849) );
  IV U2934 ( .A(n2853), .Z(n3043) );
  XNOR U2935 ( .A(n2850), .B(n3044), .Z(n2853) );
  AND U2936 ( .A(n42), .B(n9621), .Z(n3044) );
  XOR U2937 ( .A(n3045), .B(n3046), .Z(n2850) );
  ANDN U2938 ( .A(n3047), .B(n3048), .Z(n3046) );
  XNOR U2939 ( .A(n3045), .B(n3049), .Z(n3047) );
  XNOR U2940 ( .A(n3050), .B(n3051), .Z(n2854) );
  ANDN U2941 ( .A(n3052), .B(n3053), .Z(n3051) );
  XNOR U2942 ( .A(n3050), .B(n3054), .Z(n3052) );
  XNOR U2943 ( .A(n2863), .B(n2855), .Z(n2873) );
  XOR U2944 ( .A(n3055), .B(n3056), .Z(n2855) );
  AND U2945 ( .A(n3057), .B(n3058), .Z(n3056) );
  XNOR U2946 ( .A(n3059), .B(n3055), .Z(n3058) );
  XOR U2947 ( .A(n2861), .B(n3060), .Z(n2863) );
  ANDN U2948 ( .A(n9621), .B(n43), .Z(n3060) );
  XOR U2949 ( .A(n3061), .B(n3062), .Z(n2861) );
  AND U2950 ( .A(n3063), .B(n3064), .Z(n3062) );
  XNOR U2951 ( .A(n3061), .B(n3065), .Z(n3064) );
  XOR U2952 ( .A(n2859), .B(n2869), .Z(n2872) );
  XOR U2953 ( .A(n3066), .B(n3067), .Z(n2859) );
  IV U2954 ( .A(n3068), .Z(n3067) );
  XOR U2955 ( .A(n3069), .B(n3070), .Z(n2869) );
  AND U2956 ( .A(n3069), .B(n3071), .Z(n3070) );
  XOR U2957 ( .A(n3072), .B(n3057), .Z(n3071) );
  XOR U2958 ( .A(n3073), .B(n3065), .Z(n3057) );
  XOR U2959 ( .A(n2880), .B(n3074), .Z(n3065) );
  IV U2960 ( .A(n2879), .Z(n3074) );
  XNOR U2961 ( .A(n2876), .B(n3075), .Z(n2879) );
  XOR U2962 ( .A(n3076), .B(n3077), .Z(n2876) );
  ANDN U2963 ( .A(n3078), .B(n3079), .Z(n3077) );
  XNOR U2964 ( .A(n3076), .B(n3080), .Z(n3078) );
  XOR U2965 ( .A(n2887), .B(n3081), .Z(n2880) );
  IV U2966 ( .A(n2886), .Z(n3081) );
  XNOR U2967 ( .A(n2883), .B(n3082), .Z(n2886) );
  XOR U2968 ( .A(n3083), .B(n3084), .Z(n2883) );
  ANDN U2969 ( .A(n3085), .B(n3086), .Z(n3084) );
  XNOR U2970 ( .A(n3083), .B(n3087), .Z(n3085) );
  XOR U2971 ( .A(n2894), .B(n3088), .Z(n2887) );
  IV U2972 ( .A(n2893), .Z(n3088) );
  XNOR U2973 ( .A(n2890), .B(n3089), .Z(n2893) );
  XOR U2974 ( .A(n3090), .B(n3091), .Z(n2890) );
  ANDN U2975 ( .A(n3092), .B(n3093), .Z(n3091) );
  XNOR U2976 ( .A(n3090), .B(n3094), .Z(n3092) );
  XOR U2977 ( .A(n2901), .B(n3095), .Z(n2894) );
  IV U2978 ( .A(n2900), .Z(n3095) );
  XNOR U2979 ( .A(n2897), .B(n3096), .Z(n2900) );
  XOR U2980 ( .A(n3097), .B(n3098), .Z(n2897) );
  ANDN U2981 ( .A(n3099), .B(n3100), .Z(n3098) );
  XNOR U2982 ( .A(n3097), .B(n3101), .Z(n3099) );
  XOR U2983 ( .A(n2908), .B(n3102), .Z(n2901) );
  IV U2984 ( .A(n2907), .Z(n3102) );
  XNOR U2985 ( .A(n2904), .B(n3103), .Z(n2907) );
  XOR U2986 ( .A(n3104), .B(n3105), .Z(n2904) );
  ANDN U2987 ( .A(n3106), .B(n3107), .Z(n3105) );
  XNOR U2988 ( .A(n3104), .B(n3108), .Z(n3106) );
  XOR U2989 ( .A(n2915), .B(n3109), .Z(n2908) );
  IV U2990 ( .A(n2914), .Z(n3109) );
  XNOR U2991 ( .A(n2911), .B(n3110), .Z(n2914) );
  XOR U2992 ( .A(n3111), .B(n3112), .Z(n2911) );
  ANDN U2993 ( .A(n3113), .B(n3114), .Z(n3112) );
  XNOR U2994 ( .A(n3111), .B(n3115), .Z(n3113) );
  XOR U2995 ( .A(n2922), .B(n3116), .Z(n2915) );
  IV U2996 ( .A(n2921), .Z(n3116) );
  XNOR U2997 ( .A(n2918), .B(n3117), .Z(n2921) );
  XOR U2998 ( .A(n3118), .B(n3119), .Z(n2918) );
  ANDN U2999 ( .A(n3120), .B(n3121), .Z(n3119) );
  XNOR U3000 ( .A(n3118), .B(n3122), .Z(n3120) );
  XOR U3001 ( .A(n2929), .B(n3123), .Z(n2922) );
  IV U3002 ( .A(n2928), .Z(n3123) );
  XNOR U3003 ( .A(n2925), .B(n3124), .Z(n2928) );
  XOR U3004 ( .A(n3125), .B(n3126), .Z(n2925) );
  ANDN U3005 ( .A(n3127), .B(n3128), .Z(n3126) );
  XNOR U3006 ( .A(n3125), .B(n3129), .Z(n3127) );
  XOR U3007 ( .A(n2936), .B(n3130), .Z(n2929) );
  IV U3008 ( .A(n2935), .Z(n3130) );
  XNOR U3009 ( .A(n2932), .B(n3131), .Z(n2935) );
  XOR U3010 ( .A(n3132), .B(n3133), .Z(n2932) );
  ANDN U3011 ( .A(n3134), .B(n3135), .Z(n3133) );
  XNOR U3012 ( .A(n3132), .B(n3136), .Z(n3134) );
  XOR U3013 ( .A(n2943), .B(n3137), .Z(n2936) );
  IV U3014 ( .A(n2942), .Z(n3137) );
  XNOR U3015 ( .A(n2939), .B(n3138), .Z(n2942) );
  XOR U3016 ( .A(n3139), .B(n3140), .Z(n2939) );
  ANDN U3017 ( .A(n3141), .B(n3142), .Z(n3140) );
  XNOR U3018 ( .A(n3139), .B(n3143), .Z(n3141) );
  XOR U3019 ( .A(n2950), .B(n3144), .Z(n2943) );
  IV U3020 ( .A(n2949), .Z(n3144) );
  XNOR U3021 ( .A(n2946), .B(n3145), .Z(n2949) );
  XOR U3022 ( .A(n3146), .B(n3147), .Z(n2946) );
  ANDN U3023 ( .A(n3148), .B(n3149), .Z(n3147) );
  XNOR U3024 ( .A(n3146), .B(n3150), .Z(n3148) );
  XOR U3025 ( .A(n2957), .B(n3151), .Z(n2950) );
  IV U3026 ( .A(n2956), .Z(n3151) );
  XNOR U3027 ( .A(n2953), .B(n3152), .Z(n2956) );
  XOR U3028 ( .A(n3153), .B(n3154), .Z(n2953) );
  ANDN U3029 ( .A(n3155), .B(n3156), .Z(n3154) );
  XNOR U3030 ( .A(n3153), .B(n3157), .Z(n3155) );
  XOR U3031 ( .A(n2964), .B(n3158), .Z(n2957) );
  IV U3032 ( .A(n2963), .Z(n3158) );
  XNOR U3033 ( .A(n2960), .B(n3159), .Z(n2963) );
  XOR U3034 ( .A(n3160), .B(n3161), .Z(n2960) );
  ANDN U3035 ( .A(n3162), .B(n3163), .Z(n3161) );
  XNOR U3036 ( .A(n3160), .B(n3164), .Z(n3162) );
  XOR U3037 ( .A(n2970), .B(n3165), .Z(n2964) );
  IV U3038 ( .A(n2969), .Z(n3165) );
  XNOR U3039 ( .A(n2966), .B(n3166), .Z(n2969) );
  XOR U3040 ( .A(n3167), .B(n3168), .Z(n2966) );
  ANDN U3041 ( .A(n3169), .B(n3170), .Z(n3168) );
  XNOR U3042 ( .A(n3167), .B(n3171), .Z(n3169) );
  XOR U3043 ( .A(n2976), .B(n3172), .Z(n2970) );
  IV U3044 ( .A(n2975), .Z(n3172) );
  XNOR U3045 ( .A(n2972), .B(n3159), .Z(n2975) );
  AND U3046 ( .A(n3593), .B(n2765), .Z(n3159) );
  XOR U3047 ( .A(n3173), .B(n3174), .Z(n2972) );
  ANDN U3048 ( .A(n3175), .B(n3176), .Z(n3174) );
  XNOR U3049 ( .A(n3173), .B(n3177), .Z(n3175) );
  XOR U3050 ( .A(n2982), .B(n3178), .Z(n2976) );
  IV U3051 ( .A(n2981), .Z(n3178) );
  XNOR U3052 ( .A(n2978), .B(n3152), .Z(n2981) );
  AND U3053 ( .A(n4046), .B(n2396), .Z(n3152) );
  XOR U3054 ( .A(n3179), .B(n3180), .Z(n2978) );
  ANDN U3055 ( .A(n3181), .B(n3182), .Z(n3180) );
  XNOR U3056 ( .A(n3179), .B(n3183), .Z(n3181) );
  XOR U3057 ( .A(n2988), .B(n3184), .Z(n2982) );
  IV U3058 ( .A(n2987), .Z(n3184) );
  XNOR U3059 ( .A(n2984), .B(n3145), .Z(n2987) );
  AND U3060 ( .A(n4525), .B(n2053), .Z(n3145) );
  XOR U3061 ( .A(n3185), .B(n3186), .Z(n2984) );
  ANDN U3062 ( .A(n3187), .B(n3188), .Z(n3186) );
  XNOR U3063 ( .A(n3185), .B(n3189), .Z(n3187) );
  XOR U3064 ( .A(n2994), .B(n3190), .Z(n2988) );
  IV U3065 ( .A(n2993), .Z(n3190) );
  XNOR U3066 ( .A(n2990), .B(n3138), .Z(n2993) );
  AND U3067 ( .A(n5030), .B(n1737), .Z(n3138) );
  XOR U3068 ( .A(n3191), .B(n3192), .Z(n2990) );
  ANDN U3069 ( .A(n3193), .B(n3194), .Z(n3192) );
  XNOR U3070 ( .A(n3191), .B(n3195), .Z(n3193) );
  XOR U3071 ( .A(n3000), .B(n3196), .Z(n2994) );
  IV U3072 ( .A(n2999), .Z(n3196) );
  XNOR U3073 ( .A(n2996), .B(n3131), .Z(n2999) );
  AND U3074 ( .A(n5561), .B(n1448), .Z(n3131) );
  XOR U3075 ( .A(n3197), .B(n3198), .Z(n2996) );
  ANDN U3076 ( .A(n3199), .B(n3200), .Z(n3198) );
  XNOR U3077 ( .A(n3197), .B(n3201), .Z(n3199) );
  XOR U3078 ( .A(n3006), .B(n3202), .Z(n3000) );
  IV U3079 ( .A(n3005), .Z(n3202) );
  XNOR U3080 ( .A(n3002), .B(n3124), .Z(n3005) );
  AND U3081 ( .A(n6118), .B(n1185), .Z(n3124) );
  XOR U3082 ( .A(n3203), .B(n3204), .Z(n3002) );
  ANDN U3083 ( .A(n3205), .B(n3206), .Z(n3204) );
  XNOR U3084 ( .A(n3203), .B(n3207), .Z(n3205) );
  XOR U3085 ( .A(n3012), .B(n3208), .Z(n3006) );
  IV U3086 ( .A(n3011), .Z(n3208) );
  XNOR U3087 ( .A(n3008), .B(n3117), .Z(n3011) );
  AND U3088 ( .A(n6688), .B(n948), .Z(n3117) );
  XOR U3089 ( .A(n3209), .B(n3210), .Z(n3008) );
  ANDN U3090 ( .A(n3211), .B(n3212), .Z(n3210) );
  XNOR U3091 ( .A(n3209), .B(n3213), .Z(n3211) );
  XOR U3092 ( .A(n3018), .B(n3214), .Z(n3012) );
  IV U3093 ( .A(n3017), .Z(n3214) );
  XNOR U3094 ( .A(n3014), .B(n3110), .Z(n3017) );
  AND U3095 ( .A(n7241), .B(n736), .Z(n3110) );
  XOR U3096 ( .A(n3215), .B(n3216), .Z(n3014) );
  ANDN U3097 ( .A(n3217), .B(n3218), .Z(n3216) );
  XNOR U3098 ( .A(n3215), .B(n3219), .Z(n3217) );
  XOR U3099 ( .A(n3024), .B(n3220), .Z(n3018) );
  IV U3100 ( .A(n3023), .Z(n3220) );
  XNOR U3101 ( .A(n3020), .B(n3103), .Z(n3023) );
  AND U3102 ( .A(n7770), .B(n552), .Z(n3103) );
  XOR U3103 ( .A(n3221), .B(n3222), .Z(n3020) );
  ANDN U3104 ( .A(n3223), .B(n3224), .Z(n3222) );
  XNOR U3105 ( .A(n3221), .B(n3225), .Z(n3223) );
  XOR U3106 ( .A(n3030), .B(n3226), .Z(n3024) );
  IV U3107 ( .A(n3029), .Z(n3226) );
  XNOR U3108 ( .A(n3026), .B(n3096), .Z(n3029) );
  AND U3109 ( .A(n8272), .B(n395), .Z(n3096) );
  XOR U3110 ( .A(n3227), .B(n3228), .Z(n3026) );
  ANDN U3111 ( .A(n3229), .B(n3230), .Z(n3228) );
  XNOR U3112 ( .A(n3227), .B(n3231), .Z(n3229) );
  XOR U3113 ( .A(n3036), .B(n3232), .Z(n3030) );
  IV U3114 ( .A(n3035), .Z(n3232) );
  XNOR U3115 ( .A(n3032), .B(n3089), .Z(n3035) );
  AND U3116 ( .A(n8748), .B(n264), .Z(n3089) );
  XOR U3117 ( .A(n3233), .B(n3234), .Z(n3032) );
  ANDN U3118 ( .A(n3235), .B(n3236), .Z(n3234) );
  XNOR U3119 ( .A(n3233), .B(n3237), .Z(n3235) );
  XOR U3120 ( .A(n3042), .B(n3238), .Z(n3036) );
  IV U3121 ( .A(n3041), .Z(n3238) );
  XNOR U3122 ( .A(n3038), .B(n3082), .Z(n3041) );
  AND U3123 ( .A(n9198), .B(n159), .Z(n3082) );
  XOR U3124 ( .A(n3239), .B(n3240), .Z(n3038) );
  ANDN U3125 ( .A(n3241), .B(n3242), .Z(n3240) );
  XNOR U3126 ( .A(n3239), .B(n3243), .Z(n3241) );
  XOR U3127 ( .A(n3049), .B(n3244), .Z(n3042) );
  IV U3128 ( .A(n3048), .Z(n3244) );
  XNOR U3129 ( .A(n3045), .B(n3075), .Z(n3048) );
  AND U3130 ( .A(n9621), .B(n80), .Z(n3075) );
  XOR U3131 ( .A(n3245), .B(n3246), .Z(n3045) );
  ANDN U3132 ( .A(n3247), .B(n3248), .Z(n3246) );
  XNOR U3133 ( .A(n3245), .B(n3249), .Z(n3247) );
  XOR U3134 ( .A(n3054), .B(n3250), .Z(n3049) );
  IV U3135 ( .A(n3053), .Z(n3250) );
  XNOR U3136 ( .A(n3050), .B(n3251), .Z(n3053) );
  AND U3137 ( .A(n42), .B(n10017), .Z(n3251) );
  XOR U3138 ( .A(n3252), .B(n3253), .Z(n3050) );
  ANDN U3139 ( .A(n3254), .B(n3255), .Z(n3253) );
  XNOR U3140 ( .A(n3252), .B(n3256), .Z(n3254) );
  XNOR U3141 ( .A(n3257), .B(n3258), .Z(n3054) );
  ANDN U3142 ( .A(n3259), .B(n3260), .Z(n3258) );
  XNOR U3143 ( .A(n3257), .B(n3261), .Z(n3259) );
  XNOR U3144 ( .A(n3063), .B(n3055), .Z(n3073) );
  XOR U3145 ( .A(n3262), .B(n3263), .Z(n3055) );
  AND U3146 ( .A(n3264), .B(n3265), .Z(n3263) );
  XNOR U3147 ( .A(n3266), .B(n3262), .Z(n3265) );
  XOR U3148 ( .A(n3061), .B(n3267), .Z(n3063) );
  ANDN U3149 ( .A(n10017), .B(n43), .Z(n3267) );
  XOR U3150 ( .A(n3268), .B(n3269), .Z(n3061) );
  AND U3151 ( .A(n3270), .B(n3271), .Z(n3269) );
  XNOR U3152 ( .A(n3268), .B(n3272), .Z(n3271) );
  XOR U3153 ( .A(n3059), .B(n3069), .Z(n3072) );
  XOR U3154 ( .A(n3273), .B(n3274), .Z(n3059) );
  IV U3155 ( .A(n3275), .Z(n3274) );
  XOR U3156 ( .A(n3276), .B(n3277), .Z(n3069) );
  AND U3157 ( .A(n3276), .B(n3278), .Z(n3277) );
  XOR U3158 ( .A(n3279), .B(n3264), .Z(n3278) );
  XOR U3159 ( .A(n3280), .B(n3272), .Z(n3264) );
  XOR U3160 ( .A(n3080), .B(n3281), .Z(n3272) );
  IV U3161 ( .A(n3079), .Z(n3281) );
  XNOR U3162 ( .A(n3076), .B(n3282), .Z(n3079) );
  XOR U3163 ( .A(n3283), .B(n3284), .Z(n3076) );
  ANDN U3164 ( .A(n3285), .B(n3286), .Z(n3284) );
  XNOR U3165 ( .A(n3283), .B(n3287), .Z(n3285) );
  XOR U3166 ( .A(n3087), .B(n3288), .Z(n3080) );
  IV U3167 ( .A(n3086), .Z(n3288) );
  XNOR U3168 ( .A(n3083), .B(n3289), .Z(n3086) );
  XOR U3169 ( .A(n3290), .B(n3291), .Z(n3083) );
  ANDN U3170 ( .A(n3292), .B(n3293), .Z(n3291) );
  XNOR U3171 ( .A(n3290), .B(n3294), .Z(n3292) );
  XOR U3172 ( .A(n3094), .B(n3295), .Z(n3087) );
  IV U3173 ( .A(n3093), .Z(n3295) );
  XNOR U3174 ( .A(n3090), .B(n3296), .Z(n3093) );
  XOR U3175 ( .A(n3297), .B(n3298), .Z(n3090) );
  ANDN U3176 ( .A(n3299), .B(n3300), .Z(n3298) );
  XNOR U3177 ( .A(n3297), .B(n3301), .Z(n3299) );
  XOR U3178 ( .A(n3101), .B(n3302), .Z(n3094) );
  IV U3179 ( .A(n3100), .Z(n3302) );
  XNOR U3180 ( .A(n3097), .B(n3303), .Z(n3100) );
  XOR U3181 ( .A(n3304), .B(n3305), .Z(n3097) );
  ANDN U3182 ( .A(n3306), .B(n3307), .Z(n3305) );
  XNOR U3183 ( .A(n3304), .B(n3308), .Z(n3306) );
  XOR U3184 ( .A(n3108), .B(n3309), .Z(n3101) );
  IV U3185 ( .A(n3107), .Z(n3309) );
  XNOR U3186 ( .A(n3104), .B(n3310), .Z(n3107) );
  XOR U3187 ( .A(n3311), .B(n3312), .Z(n3104) );
  ANDN U3188 ( .A(n3313), .B(n3314), .Z(n3312) );
  XNOR U3189 ( .A(n3311), .B(n3315), .Z(n3313) );
  XOR U3190 ( .A(n3115), .B(n3316), .Z(n3108) );
  IV U3191 ( .A(n3114), .Z(n3316) );
  XNOR U3192 ( .A(n3111), .B(n3317), .Z(n3114) );
  XOR U3193 ( .A(n3318), .B(n3319), .Z(n3111) );
  ANDN U3194 ( .A(n3320), .B(n3321), .Z(n3319) );
  XNOR U3195 ( .A(n3318), .B(n3322), .Z(n3320) );
  XOR U3196 ( .A(n3122), .B(n3323), .Z(n3115) );
  IV U3197 ( .A(n3121), .Z(n3323) );
  XNOR U3198 ( .A(n3118), .B(n3324), .Z(n3121) );
  XOR U3199 ( .A(n3325), .B(n3326), .Z(n3118) );
  ANDN U3200 ( .A(n3327), .B(n3328), .Z(n3326) );
  XNOR U3201 ( .A(n3325), .B(n3329), .Z(n3327) );
  XOR U3202 ( .A(n3129), .B(n3330), .Z(n3122) );
  IV U3203 ( .A(n3128), .Z(n3330) );
  XNOR U3204 ( .A(n3125), .B(n3331), .Z(n3128) );
  XOR U3205 ( .A(n3332), .B(n3333), .Z(n3125) );
  ANDN U3206 ( .A(n3334), .B(n3335), .Z(n3333) );
  XNOR U3207 ( .A(n3332), .B(n3336), .Z(n3334) );
  XOR U3208 ( .A(n3136), .B(n3337), .Z(n3129) );
  IV U3209 ( .A(n3135), .Z(n3337) );
  XNOR U3210 ( .A(n3132), .B(n3338), .Z(n3135) );
  XOR U3211 ( .A(n3339), .B(n3340), .Z(n3132) );
  ANDN U3212 ( .A(n3341), .B(n3342), .Z(n3340) );
  XNOR U3213 ( .A(n3339), .B(n3343), .Z(n3341) );
  XOR U3214 ( .A(n3143), .B(n3344), .Z(n3136) );
  IV U3215 ( .A(n3142), .Z(n3344) );
  XNOR U3216 ( .A(n3139), .B(n3345), .Z(n3142) );
  XOR U3217 ( .A(n3346), .B(n3347), .Z(n3139) );
  ANDN U3218 ( .A(n3348), .B(n3349), .Z(n3347) );
  XNOR U3219 ( .A(n3346), .B(n3350), .Z(n3348) );
  XOR U3220 ( .A(n3150), .B(n3351), .Z(n3143) );
  IV U3221 ( .A(n3149), .Z(n3351) );
  XNOR U3222 ( .A(n3146), .B(n3352), .Z(n3149) );
  XOR U3223 ( .A(n3353), .B(n3354), .Z(n3146) );
  ANDN U3224 ( .A(n3355), .B(n3356), .Z(n3354) );
  XNOR U3225 ( .A(n3353), .B(n3357), .Z(n3355) );
  XOR U3226 ( .A(n3157), .B(n3358), .Z(n3150) );
  IV U3227 ( .A(n3156), .Z(n3358) );
  XNOR U3228 ( .A(n3153), .B(n3359), .Z(n3156) );
  XOR U3229 ( .A(n3360), .B(n3361), .Z(n3153) );
  ANDN U3230 ( .A(n3362), .B(n3363), .Z(n3361) );
  XNOR U3231 ( .A(n3360), .B(n3364), .Z(n3362) );
  XOR U3232 ( .A(n3164), .B(n3365), .Z(n3157) );
  IV U3233 ( .A(n3163), .Z(n3365) );
  XNOR U3234 ( .A(n3160), .B(n3366), .Z(n3163) );
  XOR U3235 ( .A(n3367), .B(n3368), .Z(n3160) );
  ANDN U3236 ( .A(n3369), .B(n3370), .Z(n3368) );
  XNOR U3237 ( .A(n3367), .B(n3371), .Z(n3369) );
  XOR U3238 ( .A(n3171), .B(n3372), .Z(n3164) );
  IV U3239 ( .A(n3170), .Z(n3372) );
  XNOR U3240 ( .A(n3167), .B(n3373), .Z(n3170) );
  XOR U3241 ( .A(n3374), .B(n3375), .Z(n3167) );
  ANDN U3242 ( .A(n3376), .B(n3377), .Z(n3375) );
  XNOR U3243 ( .A(n3374), .B(n3378), .Z(n3376) );
  XOR U3244 ( .A(n3177), .B(n3379), .Z(n3171) );
  IV U3245 ( .A(n3176), .Z(n3379) );
  XNOR U3246 ( .A(n3173), .B(n3373), .Z(n3176) );
  AND U3247 ( .A(n3593), .B(n3166), .Z(n3373) );
  XOR U3248 ( .A(n3380), .B(n3381), .Z(n3173) );
  ANDN U3249 ( .A(n3382), .B(n3383), .Z(n3381) );
  XNOR U3250 ( .A(n3380), .B(n3384), .Z(n3382) );
  XOR U3251 ( .A(n3183), .B(n3385), .Z(n3177) );
  IV U3252 ( .A(n3182), .Z(n3385) );
  XNOR U3253 ( .A(n3179), .B(n3366), .Z(n3182) );
  AND U3254 ( .A(n4046), .B(n2765), .Z(n3366) );
  XOR U3255 ( .A(n3386), .B(n3387), .Z(n3179) );
  ANDN U3256 ( .A(n3388), .B(n3389), .Z(n3387) );
  XNOR U3257 ( .A(n3386), .B(n3390), .Z(n3388) );
  XOR U3258 ( .A(n3189), .B(n3391), .Z(n3183) );
  IV U3259 ( .A(n3188), .Z(n3391) );
  XNOR U3260 ( .A(n3185), .B(n3359), .Z(n3188) );
  AND U3261 ( .A(n4525), .B(n2396), .Z(n3359) );
  XOR U3262 ( .A(n3392), .B(n3393), .Z(n3185) );
  ANDN U3263 ( .A(n3394), .B(n3395), .Z(n3393) );
  XNOR U3264 ( .A(n3392), .B(n3396), .Z(n3394) );
  XOR U3265 ( .A(n3195), .B(n3397), .Z(n3189) );
  IV U3266 ( .A(n3194), .Z(n3397) );
  XNOR U3267 ( .A(n3191), .B(n3352), .Z(n3194) );
  AND U3268 ( .A(n5030), .B(n2053), .Z(n3352) );
  XOR U3269 ( .A(n3398), .B(n3399), .Z(n3191) );
  ANDN U3270 ( .A(n3400), .B(n3401), .Z(n3399) );
  XNOR U3271 ( .A(n3398), .B(n3402), .Z(n3400) );
  XOR U3272 ( .A(n3201), .B(n3403), .Z(n3195) );
  IV U3273 ( .A(n3200), .Z(n3403) );
  XNOR U3274 ( .A(n3197), .B(n3345), .Z(n3200) );
  AND U3275 ( .A(n5561), .B(n1737), .Z(n3345) );
  XOR U3276 ( .A(n3404), .B(n3405), .Z(n3197) );
  ANDN U3277 ( .A(n3406), .B(n3407), .Z(n3405) );
  XNOR U3278 ( .A(n3404), .B(n3408), .Z(n3406) );
  XOR U3279 ( .A(n3207), .B(n3409), .Z(n3201) );
  IV U3280 ( .A(n3206), .Z(n3409) );
  XNOR U3281 ( .A(n3203), .B(n3338), .Z(n3206) );
  AND U3282 ( .A(n6118), .B(n1448), .Z(n3338) );
  XOR U3283 ( .A(n3410), .B(n3411), .Z(n3203) );
  ANDN U3284 ( .A(n3412), .B(n3413), .Z(n3411) );
  XNOR U3285 ( .A(n3410), .B(n3414), .Z(n3412) );
  XOR U3286 ( .A(n3213), .B(n3415), .Z(n3207) );
  IV U3287 ( .A(n3212), .Z(n3415) );
  XNOR U3288 ( .A(n3209), .B(n3331), .Z(n3212) );
  AND U3289 ( .A(n6688), .B(n1185), .Z(n3331) );
  XOR U3290 ( .A(n3416), .B(n3417), .Z(n3209) );
  ANDN U3291 ( .A(n3418), .B(n3419), .Z(n3417) );
  XNOR U3292 ( .A(n3416), .B(n3420), .Z(n3418) );
  XOR U3293 ( .A(n3219), .B(n3421), .Z(n3213) );
  IV U3294 ( .A(n3218), .Z(n3421) );
  XNOR U3295 ( .A(n3215), .B(n3324), .Z(n3218) );
  AND U3296 ( .A(n7241), .B(n948), .Z(n3324) );
  XOR U3297 ( .A(n3422), .B(n3423), .Z(n3215) );
  ANDN U3298 ( .A(n3424), .B(n3425), .Z(n3423) );
  XNOR U3299 ( .A(n3422), .B(n3426), .Z(n3424) );
  XOR U3300 ( .A(n3225), .B(n3427), .Z(n3219) );
  IV U3301 ( .A(n3224), .Z(n3427) );
  XNOR U3302 ( .A(n3221), .B(n3317), .Z(n3224) );
  AND U3303 ( .A(n7770), .B(n736), .Z(n3317) );
  XOR U3304 ( .A(n3428), .B(n3429), .Z(n3221) );
  ANDN U3305 ( .A(n3430), .B(n3431), .Z(n3429) );
  XNOR U3306 ( .A(n3428), .B(n3432), .Z(n3430) );
  XOR U3307 ( .A(n3231), .B(n3433), .Z(n3225) );
  IV U3308 ( .A(n3230), .Z(n3433) );
  XNOR U3309 ( .A(n3227), .B(n3310), .Z(n3230) );
  AND U3310 ( .A(n8272), .B(n552), .Z(n3310) );
  XOR U3311 ( .A(n3434), .B(n3435), .Z(n3227) );
  ANDN U3312 ( .A(n3436), .B(n3437), .Z(n3435) );
  XNOR U3313 ( .A(n3434), .B(n3438), .Z(n3436) );
  XOR U3314 ( .A(n3237), .B(n3439), .Z(n3231) );
  IV U3315 ( .A(n3236), .Z(n3439) );
  XNOR U3316 ( .A(n3233), .B(n3303), .Z(n3236) );
  AND U3317 ( .A(n8748), .B(n395), .Z(n3303) );
  XOR U3318 ( .A(n3440), .B(n3441), .Z(n3233) );
  ANDN U3319 ( .A(n3442), .B(n3443), .Z(n3441) );
  XNOR U3320 ( .A(n3440), .B(n3444), .Z(n3442) );
  XOR U3321 ( .A(n3243), .B(n3445), .Z(n3237) );
  IV U3322 ( .A(n3242), .Z(n3445) );
  XNOR U3323 ( .A(n3239), .B(n3296), .Z(n3242) );
  AND U3324 ( .A(n9198), .B(n264), .Z(n3296) );
  XOR U3325 ( .A(n3446), .B(n3447), .Z(n3239) );
  ANDN U3326 ( .A(n3448), .B(n3449), .Z(n3447) );
  XNOR U3327 ( .A(n3446), .B(n3450), .Z(n3448) );
  XOR U3328 ( .A(n3249), .B(n3451), .Z(n3243) );
  IV U3329 ( .A(n3248), .Z(n3451) );
  XNOR U3330 ( .A(n3245), .B(n3289), .Z(n3248) );
  AND U3331 ( .A(n9621), .B(n159), .Z(n3289) );
  XOR U3332 ( .A(n3452), .B(n3453), .Z(n3245) );
  ANDN U3333 ( .A(n3454), .B(n3455), .Z(n3453) );
  XNOR U3334 ( .A(n3452), .B(n3456), .Z(n3454) );
  XOR U3335 ( .A(n3256), .B(n3457), .Z(n3249) );
  IV U3336 ( .A(n3255), .Z(n3457) );
  XNOR U3337 ( .A(n3252), .B(n3282), .Z(n3255) );
  AND U3338 ( .A(n10017), .B(n80), .Z(n3282) );
  XOR U3339 ( .A(n3458), .B(n3459), .Z(n3252) );
  ANDN U3340 ( .A(n3460), .B(n3461), .Z(n3459) );
  XNOR U3341 ( .A(n3458), .B(n3462), .Z(n3460) );
  XOR U3342 ( .A(n3261), .B(n3463), .Z(n3256) );
  IV U3343 ( .A(n3260), .Z(n3463) );
  XNOR U3344 ( .A(n3257), .B(n3464), .Z(n3260) );
  AND U3345 ( .A(n42), .B(n10387), .Z(n3464) );
  XOR U3346 ( .A(n3465), .B(n3466), .Z(n3257) );
  ANDN U3347 ( .A(n3467), .B(n3468), .Z(n3466) );
  XNOR U3348 ( .A(n3465), .B(n3469), .Z(n3467) );
  XNOR U3349 ( .A(n3470), .B(n3471), .Z(n3261) );
  ANDN U3350 ( .A(n3472), .B(n3473), .Z(n3471) );
  XNOR U3351 ( .A(n3470), .B(n3474), .Z(n3472) );
  XNOR U3352 ( .A(n3270), .B(n3262), .Z(n3280) );
  XOR U3353 ( .A(n3475), .B(n3476), .Z(n3262) );
  AND U3354 ( .A(n3477), .B(n3478), .Z(n3476) );
  XNOR U3355 ( .A(n3479), .B(n3475), .Z(n3478) );
  XOR U3356 ( .A(n3268), .B(n3480), .Z(n3270) );
  ANDN U3357 ( .A(n10387), .B(n43), .Z(n3480) );
  XOR U3358 ( .A(n3481), .B(n3482), .Z(n3268) );
  AND U3359 ( .A(n3483), .B(n3484), .Z(n3482) );
  XNOR U3360 ( .A(n3481), .B(n3485), .Z(n3484) );
  XOR U3361 ( .A(n3266), .B(n3276), .Z(n3279) );
  XOR U3362 ( .A(n3486), .B(n3487), .Z(n3266) );
  IV U3363 ( .A(n3488), .Z(n3487) );
  XOR U3364 ( .A(n3489), .B(n3490), .Z(n3276) );
  AND U3365 ( .A(n3489), .B(n3491), .Z(n3490) );
  XOR U3366 ( .A(n3492), .B(n3477), .Z(n3491) );
  XOR U3367 ( .A(n3493), .B(n3485), .Z(n3477) );
  XOR U3368 ( .A(n3287), .B(n3494), .Z(n3485) );
  IV U3369 ( .A(n3286), .Z(n3494) );
  XNOR U3370 ( .A(n3283), .B(n3495), .Z(n3286) );
  XOR U3371 ( .A(n3496), .B(n3497), .Z(n3283) );
  ANDN U3372 ( .A(n3498), .B(n3499), .Z(n3497) );
  XNOR U3373 ( .A(n3496), .B(n3500), .Z(n3498) );
  XOR U3374 ( .A(n3294), .B(n3501), .Z(n3287) );
  IV U3375 ( .A(n3293), .Z(n3501) );
  XNOR U3376 ( .A(n3290), .B(n3502), .Z(n3293) );
  XOR U3377 ( .A(n3503), .B(n3504), .Z(n3290) );
  ANDN U3378 ( .A(n3505), .B(n3506), .Z(n3504) );
  XNOR U3379 ( .A(n3503), .B(n3507), .Z(n3505) );
  XOR U3380 ( .A(n3301), .B(n3508), .Z(n3294) );
  IV U3381 ( .A(n3300), .Z(n3508) );
  XNOR U3382 ( .A(n3297), .B(n3509), .Z(n3300) );
  XOR U3383 ( .A(n3510), .B(n3511), .Z(n3297) );
  ANDN U3384 ( .A(n3512), .B(n3513), .Z(n3511) );
  XNOR U3385 ( .A(n3510), .B(n3514), .Z(n3512) );
  XOR U3386 ( .A(n3308), .B(n3515), .Z(n3301) );
  IV U3387 ( .A(n3307), .Z(n3515) );
  XNOR U3388 ( .A(n3304), .B(n3516), .Z(n3307) );
  XOR U3389 ( .A(n3517), .B(n3518), .Z(n3304) );
  ANDN U3390 ( .A(n3519), .B(n3520), .Z(n3518) );
  XNOR U3391 ( .A(n3517), .B(n3521), .Z(n3519) );
  XOR U3392 ( .A(n3315), .B(n3522), .Z(n3308) );
  IV U3393 ( .A(n3314), .Z(n3522) );
  XNOR U3394 ( .A(n3311), .B(n3523), .Z(n3314) );
  XOR U3395 ( .A(n3524), .B(n3525), .Z(n3311) );
  ANDN U3396 ( .A(n3526), .B(n3527), .Z(n3525) );
  XNOR U3397 ( .A(n3524), .B(n3528), .Z(n3526) );
  XOR U3398 ( .A(n3322), .B(n3529), .Z(n3315) );
  IV U3399 ( .A(n3321), .Z(n3529) );
  XNOR U3400 ( .A(n3318), .B(n3530), .Z(n3321) );
  XOR U3401 ( .A(n3531), .B(n3532), .Z(n3318) );
  ANDN U3402 ( .A(n3533), .B(n3534), .Z(n3532) );
  XNOR U3403 ( .A(n3531), .B(n3535), .Z(n3533) );
  XOR U3404 ( .A(n3329), .B(n3536), .Z(n3322) );
  IV U3405 ( .A(n3328), .Z(n3536) );
  XNOR U3406 ( .A(n3325), .B(n3537), .Z(n3328) );
  XOR U3407 ( .A(n3538), .B(n3539), .Z(n3325) );
  ANDN U3408 ( .A(n3540), .B(n3541), .Z(n3539) );
  XNOR U3409 ( .A(n3538), .B(n3542), .Z(n3540) );
  XOR U3410 ( .A(n3336), .B(n3543), .Z(n3329) );
  IV U3411 ( .A(n3335), .Z(n3543) );
  XNOR U3412 ( .A(n3332), .B(n3544), .Z(n3335) );
  XOR U3413 ( .A(n3545), .B(n3546), .Z(n3332) );
  ANDN U3414 ( .A(n3547), .B(n3548), .Z(n3546) );
  XNOR U3415 ( .A(n3545), .B(n3549), .Z(n3547) );
  XOR U3416 ( .A(n3343), .B(n3550), .Z(n3336) );
  IV U3417 ( .A(n3342), .Z(n3550) );
  XNOR U3418 ( .A(n3339), .B(n3551), .Z(n3342) );
  XOR U3419 ( .A(n3552), .B(n3553), .Z(n3339) );
  ANDN U3420 ( .A(n3554), .B(n3555), .Z(n3553) );
  XNOR U3421 ( .A(n3552), .B(n3556), .Z(n3554) );
  XOR U3422 ( .A(n3350), .B(n3557), .Z(n3343) );
  IV U3423 ( .A(n3349), .Z(n3557) );
  XNOR U3424 ( .A(n3346), .B(n3558), .Z(n3349) );
  XOR U3425 ( .A(n3559), .B(n3560), .Z(n3346) );
  ANDN U3426 ( .A(n3561), .B(n3562), .Z(n3560) );
  XNOR U3427 ( .A(n3559), .B(n3563), .Z(n3561) );
  XOR U3428 ( .A(n3357), .B(n3564), .Z(n3350) );
  IV U3429 ( .A(n3356), .Z(n3564) );
  XNOR U3430 ( .A(n3353), .B(n3565), .Z(n3356) );
  XOR U3431 ( .A(n3566), .B(n3567), .Z(n3353) );
  ANDN U3432 ( .A(n3568), .B(n3569), .Z(n3567) );
  XNOR U3433 ( .A(n3566), .B(n3570), .Z(n3568) );
  XOR U3434 ( .A(n3364), .B(n3571), .Z(n3357) );
  IV U3435 ( .A(n3363), .Z(n3571) );
  XNOR U3436 ( .A(n3360), .B(n3572), .Z(n3363) );
  XOR U3437 ( .A(n3573), .B(n3574), .Z(n3360) );
  ANDN U3438 ( .A(n3575), .B(n3576), .Z(n3574) );
  XNOR U3439 ( .A(n3573), .B(n3577), .Z(n3575) );
  XOR U3440 ( .A(n3371), .B(n3578), .Z(n3364) );
  IV U3441 ( .A(n3370), .Z(n3578) );
  XNOR U3442 ( .A(n3367), .B(n3579), .Z(n3370) );
  XOR U3443 ( .A(n3580), .B(n3581), .Z(n3367) );
  ANDN U3444 ( .A(n3582), .B(n3583), .Z(n3581) );
  XNOR U3445 ( .A(n3580), .B(n3584), .Z(n3582) );
  XOR U3446 ( .A(n3378), .B(n3585), .Z(n3371) );
  IV U3447 ( .A(n3377), .Z(n3585) );
  XNOR U3448 ( .A(n3374), .B(n3586), .Z(n3377) );
  XOR U3449 ( .A(n3587), .B(n3588), .Z(n3374) );
  ANDN U3450 ( .A(n3589), .B(n3590), .Z(n3588) );
  XNOR U3451 ( .A(n3587), .B(n3591), .Z(n3589) );
  XOR U3452 ( .A(n3384), .B(n3592), .Z(n3378) );
  IV U3453 ( .A(n3383), .Z(n3592) );
  XNOR U3454 ( .A(n3380), .B(n3593), .Z(n3383) );
  XOR U3455 ( .A(n3594), .B(n3595), .Z(n3380) );
  ANDN U3456 ( .A(n3596), .B(n3597), .Z(n3595) );
  XNOR U3457 ( .A(n3594), .B(n3598), .Z(n3596) );
  XOR U3458 ( .A(n3390), .B(n3599), .Z(n3384) );
  IV U3459 ( .A(n3389), .Z(n3599) );
  XNOR U3460 ( .A(n3386), .B(n3586), .Z(n3389) );
  AND U3461 ( .A(n4046), .B(n3166), .Z(n3586) );
  XOR U3462 ( .A(n3600), .B(n3601), .Z(n3386) );
  ANDN U3463 ( .A(n3602), .B(n3603), .Z(n3601) );
  XNOR U3464 ( .A(n3600), .B(n3604), .Z(n3602) );
  XOR U3465 ( .A(n3396), .B(n3605), .Z(n3390) );
  IV U3466 ( .A(n3395), .Z(n3605) );
  XNOR U3467 ( .A(n3392), .B(n3579), .Z(n3395) );
  AND U3468 ( .A(n4525), .B(n2765), .Z(n3579) );
  XOR U3469 ( .A(n3606), .B(n3607), .Z(n3392) );
  ANDN U3470 ( .A(n3608), .B(n3609), .Z(n3607) );
  XNOR U3471 ( .A(n3606), .B(n3610), .Z(n3608) );
  XOR U3472 ( .A(n3402), .B(n3611), .Z(n3396) );
  IV U3473 ( .A(n3401), .Z(n3611) );
  XNOR U3474 ( .A(n3398), .B(n3572), .Z(n3401) );
  AND U3475 ( .A(n5030), .B(n2396), .Z(n3572) );
  XOR U3476 ( .A(n3612), .B(n3613), .Z(n3398) );
  ANDN U3477 ( .A(n3614), .B(n3615), .Z(n3613) );
  XNOR U3478 ( .A(n3612), .B(n3616), .Z(n3614) );
  XOR U3479 ( .A(n3408), .B(n3617), .Z(n3402) );
  IV U3480 ( .A(n3407), .Z(n3617) );
  XNOR U3481 ( .A(n3404), .B(n3565), .Z(n3407) );
  AND U3482 ( .A(n5561), .B(n2053), .Z(n3565) );
  XOR U3483 ( .A(n3618), .B(n3619), .Z(n3404) );
  ANDN U3484 ( .A(n3620), .B(n3621), .Z(n3619) );
  XNOR U3485 ( .A(n3618), .B(n3622), .Z(n3620) );
  XOR U3486 ( .A(n3414), .B(n3623), .Z(n3408) );
  IV U3487 ( .A(n3413), .Z(n3623) );
  XNOR U3488 ( .A(n3410), .B(n3558), .Z(n3413) );
  AND U3489 ( .A(n6118), .B(n1737), .Z(n3558) );
  XOR U3490 ( .A(n3624), .B(n3625), .Z(n3410) );
  ANDN U3491 ( .A(n3626), .B(n3627), .Z(n3625) );
  XNOR U3492 ( .A(n3624), .B(n3628), .Z(n3626) );
  XOR U3493 ( .A(n3420), .B(n3629), .Z(n3414) );
  IV U3494 ( .A(n3419), .Z(n3629) );
  XNOR U3495 ( .A(n3416), .B(n3551), .Z(n3419) );
  AND U3496 ( .A(n6688), .B(n1448), .Z(n3551) );
  XOR U3497 ( .A(n3630), .B(n3631), .Z(n3416) );
  ANDN U3498 ( .A(n3632), .B(n3633), .Z(n3631) );
  XNOR U3499 ( .A(n3630), .B(n3634), .Z(n3632) );
  XOR U3500 ( .A(n3426), .B(n3635), .Z(n3420) );
  IV U3501 ( .A(n3425), .Z(n3635) );
  XNOR U3502 ( .A(n3422), .B(n3544), .Z(n3425) );
  AND U3503 ( .A(n7241), .B(n1185), .Z(n3544) );
  XOR U3504 ( .A(n3636), .B(n3637), .Z(n3422) );
  ANDN U3505 ( .A(n3638), .B(n3639), .Z(n3637) );
  XNOR U3506 ( .A(n3636), .B(n3640), .Z(n3638) );
  XOR U3507 ( .A(n3432), .B(n3641), .Z(n3426) );
  IV U3508 ( .A(n3431), .Z(n3641) );
  XNOR U3509 ( .A(n3428), .B(n3537), .Z(n3431) );
  AND U3510 ( .A(n7770), .B(n948), .Z(n3537) );
  XOR U3511 ( .A(n3642), .B(n3643), .Z(n3428) );
  ANDN U3512 ( .A(n3644), .B(n3645), .Z(n3643) );
  XNOR U3513 ( .A(n3642), .B(n3646), .Z(n3644) );
  XOR U3514 ( .A(n3438), .B(n3647), .Z(n3432) );
  IV U3515 ( .A(n3437), .Z(n3647) );
  XNOR U3516 ( .A(n3434), .B(n3530), .Z(n3437) );
  AND U3517 ( .A(n8272), .B(n736), .Z(n3530) );
  XOR U3518 ( .A(n3648), .B(n3649), .Z(n3434) );
  ANDN U3519 ( .A(n3650), .B(n3651), .Z(n3649) );
  XNOR U3520 ( .A(n3648), .B(n3652), .Z(n3650) );
  XOR U3521 ( .A(n3444), .B(n3653), .Z(n3438) );
  IV U3522 ( .A(n3443), .Z(n3653) );
  XNOR U3523 ( .A(n3440), .B(n3523), .Z(n3443) );
  AND U3524 ( .A(n8748), .B(n552), .Z(n3523) );
  XOR U3525 ( .A(n3654), .B(n3655), .Z(n3440) );
  ANDN U3526 ( .A(n3656), .B(n3657), .Z(n3655) );
  XNOR U3527 ( .A(n3654), .B(n3658), .Z(n3656) );
  XOR U3528 ( .A(n3450), .B(n3659), .Z(n3444) );
  IV U3529 ( .A(n3449), .Z(n3659) );
  XNOR U3530 ( .A(n3446), .B(n3516), .Z(n3449) );
  AND U3531 ( .A(n9198), .B(n395), .Z(n3516) );
  XOR U3532 ( .A(n3660), .B(n3661), .Z(n3446) );
  ANDN U3533 ( .A(n3662), .B(n3663), .Z(n3661) );
  XNOR U3534 ( .A(n3660), .B(n3664), .Z(n3662) );
  XOR U3535 ( .A(n3456), .B(n3665), .Z(n3450) );
  IV U3536 ( .A(n3455), .Z(n3665) );
  XNOR U3537 ( .A(n3452), .B(n3509), .Z(n3455) );
  AND U3538 ( .A(n9621), .B(n264), .Z(n3509) );
  XOR U3539 ( .A(n3666), .B(n3667), .Z(n3452) );
  ANDN U3540 ( .A(n3668), .B(n3669), .Z(n3667) );
  XNOR U3541 ( .A(n3666), .B(n3670), .Z(n3668) );
  XOR U3542 ( .A(n3462), .B(n3671), .Z(n3456) );
  IV U3543 ( .A(n3461), .Z(n3671) );
  XNOR U3544 ( .A(n3458), .B(n3502), .Z(n3461) );
  AND U3545 ( .A(n10017), .B(n159), .Z(n3502) );
  XOR U3546 ( .A(n3672), .B(n3673), .Z(n3458) );
  ANDN U3547 ( .A(n3674), .B(n3675), .Z(n3673) );
  XNOR U3548 ( .A(n3672), .B(n3676), .Z(n3674) );
  XOR U3549 ( .A(n3469), .B(n3677), .Z(n3462) );
  IV U3550 ( .A(n3468), .Z(n3677) );
  XNOR U3551 ( .A(n3465), .B(n3495), .Z(n3468) );
  AND U3552 ( .A(n10387), .B(n80), .Z(n3495) );
  XOR U3553 ( .A(n3678), .B(n3679), .Z(n3465) );
  ANDN U3554 ( .A(n3680), .B(n3681), .Z(n3679) );
  XNOR U3555 ( .A(n3678), .B(n3682), .Z(n3680) );
  XOR U3556 ( .A(n3474), .B(n3683), .Z(n3469) );
  IV U3557 ( .A(n3473), .Z(n3683) );
  XNOR U3558 ( .A(n3470), .B(n3684), .Z(n3473) );
  AND U3559 ( .A(n42), .B(n10731), .Z(n3684) );
  XOR U3560 ( .A(n3685), .B(n3686), .Z(n3470) );
  ANDN U3561 ( .A(n3687), .B(n3688), .Z(n3686) );
  XNOR U3562 ( .A(n3685), .B(n3689), .Z(n3687) );
  XNOR U3563 ( .A(n3690), .B(n3691), .Z(n3474) );
  ANDN U3564 ( .A(n3692), .B(n3693), .Z(n3691) );
  XNOR U3565 ( .A(n3690), .B(n3694), .Z(n3692) );
  XNOR U3566 ( .A(n3483), .B(n3475), .Z(n3493) );
  XOR U3567 ( .A(n3695), .B(n3696), .Z(n3475) );
  AND U3568 ( .A(n3697), .B(n3698), .Z(n3696) );
  XNOR U3569 ( .A(n3699), .B(n3695), .Z(n3698) );
  XOR U3570 ( .A(n3481), .B(n3700), .Z(n3483) );
  ANDN U3571 ( .A(n10731), .B(n43), .Z(n3700) );
  XOR U3572 ( .A(n3701), .B(n3702), .Z(n3481) );
  AND U3573 ( .A(n3703), .B(n3704), .Z(n3702) );
  XNOR U3574 ( .A(n3701), .B(n3705), .Z(n3704) );
  XOR U3575 ( .A(n3479), .B(n3489), .Z(n3492) );
  XOR U3576 ( .A(n3706), .B(n3707), .Z(n3479) );
  IV U3577 ( .A(n3708), .Z(n3707) );
  XOR U3578 ( .A(n3709), .B(n3710), .Z(n3489) );
  AND U3579 ( .A(n3709), .B(n3711), .Z(n3710) );
  XOR U3580 ( .A(n3712), .B(n3697), .Z(n3711) );
  XOR U3581 ( .A(n3713), .B(n3705), .Z(n3697) );
  XOR U3582 ( .A(n3500), .B(n3714), .Z(n3705) );
  IV U3583 ( .A(n3499), .Z(n3714) );
  XNOR U3584 ( .A(n3496), .B(n3715), .Z(n3499) );
  XOR U3585 ( .A(n3716), .B(n3717), .Z(n3496) );
  ANDN U3586 ( .A(n3718), .B(n3719), .Z(n3717) );
  XNOR U3587 ( .A(n3716), .B(n3720), .Z(n3718) );
  XOR U3588 ( .A(n3507), .B(n3721), .Z(n3500) );
  IV U3589 ( .A(n3506), .Z(n3721) );
  XNOR U3590 ( .A(n3503), .B(n3722), .Z(n3506) );
  XOR U3591 ( .A(n3723), .B(n3724), .Z(n3503) );
  ANDN U3592 ( .A(n3725), .B(n3726), .Z(n3724) );
  XNOR U3593 ( .A(n3723), .B(n3727), .Z(n3725) );
  XOR U3594 ( .A(n3514), .B(n3728), .Z(n3507) );
  IV U3595 ( .A(n3513), .Z(n3728) );
  XNOR U3596 ( .A(n3510), .B(n3729), .Z(n3513) );
  XOR U3597 ( .A(n3730), .B(n3731), .Z(n3510) );
  ANDN U3598 ( .A(n3732), .B(n3733), .Z(n3731) );
  XNOR U3599 ( .A(n3730), .B(n3734), .Z(n3732) );
  XOR U3600 ( .A(n3521), .B(n3735), .Z(n3514) );
  IV U3601 ( .A(n3520), .Z(n3735) );
  XNOR U3602 ( .A(n3517), .B(n3736), .Z(n3520) );
  XOR U3603 ( .A(n3737), .B(n3738), .Z(n3517) );
  ANDN U3604 ( .A(n3739), .B(n3740), .Z(n3738) );
  XNOR U3605 ( .A(n3737), .B(n3741), .Z(n3739) );
  XOR U3606 ( .A(n3528), .B(n3742), .Z(n3521) );
  IV U3607 ( .A(n3527), .Z(n3742) );
  XNOR U3608 ( .A(n3524), .B(n3743), .Z(n3527) );
  XOR U3609 ( .A(n3744), .B(n3745), .Z(n3524) );
  ANDN U3610 ( .A(n3746), .B(n3747), .Z(n3745) );
  XNOR U3611 ( .A(n3744), .B(n3748), .Z(n3746) );
  XOR U3612 ( .A(n3535), .B(n3749), .Z(n3528) );
  IV U3613 ( .A(n3534), .Z(n3749) );
  XNOR U3614 ( .A(n3531), .B(n3750), .Z(n3534) );
  XOR U3615 ( .A(n3751), .B(n3752), .Z(n3531) );
  ANDN U3616 ( .A(n3753), .B(n3754), .Z(n3752) );
  XNOR U3617 ( .A(n3751), .B(n3755), .Z(n3753) );
  XOR U3618 ( .A(n3542), .B(n3756), .Z(n3535) );
  IV U3619 ( .A(n3541), .Z(n3756) );
  XNOR U3620 ( .A(n3538), .B(n3757), .Z(n3541) );
  XOR U3621 ( .A(n3758), .B(n3759), .Z(n3538) );
  ANDN U3622 ( .A(n3760), .B(n3761), .Z(n3759) );
  XNOR U3623 ( .A(n3758), .B(n3762), .Z(n3760) );
  XOR U3624 ( .A(n3549), .B(n3763), .Z(n3542) );
  IV U3625 ( .A(n3548), .Z(n3763) );
  XNOR U3626 ( .A(n3545), .B(n3764), .Z(n3548) );
  XOR U3627 ( .A(n3765), .B(n3766), .Z(n3545) );
  ANDN U3628 ( .A(n3767), .B(n3768), .Z(n3766) );
  XNOR U3629 ( .A(n3765), .B(n3769), .Z(n3767) );
  XOR U3630 ( .A(n3556), .B(n3770), .Z(n3549) );
  IV U3631 ( .A(n3555), .Z(n3770) );
  XNOR U3632 ( .A(n3552), .B(n3771), .Z(n3555) );
  XOR U3633 ( .A(n3772), .B(n3773), .Z(n3552) );
  ANDN U3634 ( .A(n3774), .B(n3775), .Z(n3773) );
  XNOR U3635 ( .A(n3772), .B(n3776), .Z(n3774) );
  XOR U3636 ( .A(n3563), .B(n3777), .Z(n3556) );
  IV U3637 ( .A(n3562), .Z(n3777) );
  XNOR U3638 ( .A(n3559), .B(n3778), .Z(n3562) );
  XOR U3639 ( .A(n3779), .B(n3780), .Z(n3559) );
  ANDN U3640 ( .A(n3781), .B(n3782), .Z(n3780) );
  XNOR U3641 ( .A(n3779), .B(n3783), .Z(n3781) );
  XOR U3642 ( .A(n3570), .B(n3784), .Z(n3563) );
  IV U3643 ( .A(n3569), .Z(n3784) );
  XNOR U3644 ( .A(n3566), .B(n3785), .Z(n3569) );
  XOR U3645 ( .A(n3786), .B(n3787), .Z(n3566) );
  ANDN U3646 ( .A(n3788), .B(n3789), .Z(n3787) );
  XNOR U3647 ( .A(n3786), .B(n3790), .Z(n3788) );
  XOR U3648 ( .A(n3577), .B(n3791), .Z(n3570) );
  IV U3649 ( .A(n3576), .Z(n3791) );
  XNOR U3650 ( .A(n3573), .B(n3792), .Z(n3576) );
  XOR U3651 ( .A(n3793), .B(n3794), .Z(n3573) );
  ANDN U3652 ( .A(n3795), .B(n3796), .Z(n3794) );
  XNOR U3653 ( .A(n3793), .B(n3797), .Z(n3795) );
  XOR U3654 ( .A(n3584), .B(n3798), .Z(n3577) );
  IV U3655 ( .A(n3583), .Z(n3798) );
  XNOR U3656 ( .A(n3580), .B(n3799), .Z(n3583) );
  XOR U3657 ( .A(n3800), .B(n3801), .Z(n3580) );
  ANDN U3658 ( .A(n3802), .B(n3803), .Z(n3801) );
  XNOR U3659 ( .A(n3800), .B(n3804), .Z(n3802) );
  XOR U3660 ( .A(n3591), .B(n3805), .Z(n3584) );
  IV U3661 ( .A(n3590), .Z(n3805) );
  XNOR U3662 ( .A(n3587), .B(n3806), .Z(n3590) );
  XOR U3663 ( .A(n3807), .B(n3808), .Z(n3587) );
  ANDN U3664 ( .A(n3809), .B(n3810), .Z(n3808) );
  XNOR U3665 ( .A(n3807), .B(n3811), .Z(n3809) );
  XOR U3666 ( .A(n3598), .B(n3812), .Z(n3591) );
  IV U3667 ( .A(n3597), .Z(n3812) );
  XNOR U3668 ( .A(n3594), .B(n3813), .Z(n3597) );
  XOR U3669 ( .A(n3814), .B(n3815), .Z(n3594) );
  ANDN U3670 ( .A(n3816), .B(n3817), .Z(n3815) );
  XNOR U3671 ( .A(n3814), .B(n3818), .Z(n3816) );
  XOR U3672 ( .A(n3604), .B(n3819), .Z(n3598) );
  IV U3673 ( .A(n3603), .Z(n3819) );
  XNOR U3674 ( .A(n3600), .B(n3813), .Z(n3603) );
  AND U3675 ( .A(n4046), .B(n3593), .Z(n3813) );
  XOR U3676 ( .A(n3820), .B(n3821), .Z(n3600) );
  ANDN U3677 ( .A(n3822), .B(n3823), .Z(n3821) );
  XNOR U3678 ( .A(n3820), .B(n3824), .Z(n3822) );
  XOR U3679 ( .A(n3610), .B(n3825), .Z(n3604) );
  IV U3680 ( .A(n3609), .Z(n3825) );
  XNOR U3681 ( .A(n3606), .B(n3806), .Z(n3609) );
  AND U3682 ( .A(n4525), .B(n3166), .Z(n3806) );
  XOR U3683 ( .A(n3826), .B(n3827), .Z(n3606) );
  ANDN U3684 ( .A(n3828), .B(n3829), .Z(n3827) );
  XNOR U3685 ( .A(n3826), .B(n3830), .Z(n3828) );
  XOR U3686 ( .A(n3616), .B(n3831), .Z(n3610) );
  IV U3687 ( .A(n3615), .Z(n3831) );
  XNOR U3688 ( .A(n3612), .B(n3799), .Z(n3615) );
  AND U3689 ( .A(n5030), .B(n2765), .Z(n3799) );
  XOR U3690 ( .A(n3832), .B(n3833), .Z(n3612) );
  ANDN U3691 ( .A(n3834), .B(n3835), .Z(n3833) );
  XNOR U3692 ( .A(n3832), .B(n3836), .Z(n3834) );
  XOR U3693 ( .A(n3622), .B(n3837), .Z(n3616) );
  IV U3694 ( .A(n3621), .Z(n3837) );
  XNOR U3695 ( .A(n3618), .B(n3792), .Z(n3621) );
  AND U3696 ( .A(n5561), .B(n2396), .Z(n3792) );
  XOR U3697 ( .A(n3838), .B(n3839), .Z(n3618) );
  ANDN U3698 ( .A(n3840), .B(n3841), .Z(n3839) );
  XNOR U3699 ( .A(n3838), .B(n3842), .Z(n3840) );
  XOR U3700 ( .A(n3628), .B(n3843), .Z(n3622) );
  IV U3701 ( .A(n3627), .Z(n3843) );
  XNOR U3702 ( .A(n3624), .B(n3785), .Z(n3627) );
  AND U3703 ( .A(n6118), .B(n2053), .Z(n3785) );
  XOR U3704 ( .A(n3844), .B(n3845), .Z(n3624) );
  ANDN U3705 ( .A(n3846), .B(n3847), .Z(n3845) );
  XNOR U3706 ( .A(n3844), .B(n3848), .Z(n3846) );
  XOR U3707 ( .A(n3634), .B(n3849), .Z(n3628) );
  IV U3708 ( .A(n3633), .Z(n3849) );
  XNOR U3709 ( .A(n3630), .B(n3778), .Z(n3633) );
  AND U3710 ( .A(n6688), .B(n1737), .Z(n3778) );
  XOR U3711 ( .A(n3850), .B(n3851), .Z(n3630) );
  ANDN U3712 ( .A(n3852), .B(n3853), .Z(n3851) );
  XNOR U3713 ( .A(n3850), .B(n3854), .Z(n3852) );
  XOR U3714 ( .A(n3640), .B(n3855), .Z(n3634) );
  IV U3715 ( .A(n3639), .Z(n3855) );
  XNOR U3716 ( .A(n3636), .B(n3771), .Z(n3639) );
  AND U3717 ( .A(n7241), .B(n1448), .Z(n3771) );
  XOR U3718 ( .A(n3856), .B(n3857), .Z(n3636) );
  ANDN U3719 ( .A(n3858), .B(n3859), .Z(n3857) );
  XNOR U3720 ( .A(n3856), .B(n3860), .Z(n3858) );
  XOR U3721 ( .A(n3646), .B(n3861), .Z(n3640) );
  IV U3722 ( .A(n3645), .Z(n3861) );
  XNOR U3723 ( .A(n3642), .B(n3764), .Z(n3645) );
  AND U3724 ( .A(n7770), .B(n1185), .Z(n3764) );
  XOR U3725 ( .A(n3862), .B(n3863), .Z(n3642) );
  ANDN U3726 ( .A(n3864), .B(n3865), .Z(n3863) );
  XNOR U3727 ( .A(n3862), .B(n3866), .Z(n3864) );
  XOR U3728 ( .A(n3652), .B(n3867), .Z(n3646) );
  IV U3729 ( .A(n3651), .Z(n3867) );
  XNOR U3730 ( .A(n3648), .B(n3757), .Z(n3651) );
  AND U3731 ( .A(n8272), .B(n948), .Z(n3757) );
  XOR U3732 ( .A(n3868), .B(n3869), .Z(n3648) );
  ANDN U3733 ( .A(n3870), .B(n3871), .Z(n3869) );
  XNOR U3734 ( .A(n3868), .B(n3872), .Z(n3870) );
  XOR U3735 ( .A(n3658), .B(n3873), .Z(n3652) );
  IV U3736 ( .A(n3657), .Z(n3873) );
  XNOR U3737 ( .A(n3654), .B(n3750), .Z(n3657) );
  AND U3738 ( .A(n8748), .B(n736), .Z(n3750) );
  XOR U3739 ( .A(n3874), .B(n3875), .Z(n3654) );
  ANDN U3740 ( .A(n3876), .B(n3877), .Z(n3875) );
  XNOR U3741 ( .A(n3874), .B(n3878), .Z(n3876) );
  XOR U3742 ( .A(n3664), .B(n3879), .Z(n3658) );
  IV U3743 ( .A(n3663), .Z(n3879) );
  XNOR U3744 ( .A(n3660), .B(n3743), .Z(n3663) );
  AND U3745 ( .A(n9198), .B(n552), .Z(n3743) );
  XOR U3746 ( .A(n3880), .B(n3881), .Z(n3660) );
  ANDN U3747 ( .A(n3882), .B(n3883), .Z(n3881) );
  XNOR U3748 ( .A(n3880), .B(n3884), .Z(n3882) );
  XOR U3749 ( .A(n3670), .B(n3885), .Z(n3664) );
  IV U3750 ( .A(n3669), .Z(n3885) );
  XNOR U3751 ( .A(n3666), .B(n3736), .Z(n3669) );
  AND U3752 ( .A(n9621), .B(n395), .Z(n3736) );
  XOR U3753 ( .A(n3886), .B(n3887), .Z(n3666) );
  ANDN U3754 ( .A(n3888), .B(n3889), .Z(n3887) );
  XNOR U3755 ( .A(n3886), .B(n3890), .Z(n3888) );
  XOR U3756 ( .A(n3676), .B(n3891), .Z(n3670) );
  IV U3757 ( .A(n3675), .Z(n3891) );
  XNOR U3758 ( .A(n3672), .B(n3729), .Z(n3675) );
  AND U3759 ( .A(n10017), .B(n264), .Z(n3729) );
  XOR U3760 ( .A(n3892), .B(n3893), .Z(n3672) );
  ANDN U3761 ( .A(n3894), .B(n3895), .Z(n3893) );
  XNOR U3762 ( .A(n3892), .B(n3896), .Z(n3894) );
  XOR U3763 ( .A(n3682), .B(n3897), .Z(n3676) );
  IV U3764 ( .A(n3681), .Z(n3897) );
  XNOR U3765 ( .A(n3678), .B(n3722), .Z(n3681) );
  AND U3766 ( .A(n10387), .B(n159), .Z(n3722) );
  XOR U3767 ( .A(n3898), .B(n3899), .Z(n3678) );
  ANDN U3768 ( .A(n3900), .B(n3901), .Z(n3899) );
  XNOR U3769 ( .A(n3898), .B(n3902), .Z(n3900) );
  XOR U3770 ( .A(n3689), .B(n3903), .Z(n3682) );
  IV U3771 ( .A(n3688), .Z(n3903) );
  XNOR U3772 ( .A(n3685), .B(n3715), .Z(n3688) );
  AND U3773 ( .A(n10731), .B(n80), .Z(n3715) );
  XOR U3774 ( .A(n3904), .B(n3905), .Z(n3685) );
  ANDN U3775 ( .A(n3906), .B(n3907), .Z(n3905) );
  XNOR U3776 ( .A(n3904), .B(n3908), .Z(n3906) );
  XOR U3777 ( .A(n3694), .B(n3909), .Z(n3689) );
  IV U3778 ( .A(n3693), .Z(n3909) );
  XNOR U3779 ( .A(n3690), .B(n3910), .Z(n3693) );
  AND U3780 ( .A(n42), .B(n11049), .Z(n3910) );
  XOR U3781 ( .A(n3911), .B(n3912), .Z(n3690) );
  ANDN U3782 ( .A(n3913), .B(n3914), .Z(n3912) );
  XNOR U3783 ( .A(n3911), .B(n3915), .Z(n3913) );
  XNOR U3784 ( .A(n3916), .B(n3917), .Z(n3694) );
  ANDN U3785 ( .A(n3918), .B(n3919), .Z(n3917) );
  XNOR U3786 ( .A(n3916), .B(n3920), .Z(n3918) );
  XNOR U3787 ( .A(n3703), .B(n3695), .Z(n3713) );
  XOR U3788 ( .A(n3921), .B(n3922), .Z(n3695) );
  AND U3789 ( .A(n3923), .B(n3924), .Z(n3922) );
  XNOR U3790 ( .A(n3925), .B(n3921), .Z(n3924) );
  XOR U3791 ( .A(n3701), .B(n3926), .Z(n3703) );
  ANDN U3792 ( .A(n11049), .B(n43), .Z(n3926) );
  XOR U3793 ( .A(n3927), .B(n3928), .Z(n3701) );
  AND U3794 ( .A(n3929), .B(n3930), .Z(n3928) );
  XNOR U3795 ( .A(n3927), .B(n3931), .Z(n3930) );
  XOR U3796 ( .A(n3699), .B(n3709), .Z(n3712) );
  XOR U3797 ( .A(n3932), .B(n3933), .Z(n3699) );
  IV U3798 ( .A(n3934), .Z(n3933) );
  XOR U3799 ( .A(n3935), .B(n3936), .Z(n3709) );
  AND U3800 ( .A(n3935), .B(n3937), .Z(n3936) );
  XOR U3801 ( .A(n3938), .B(n3923), .Z(n3937) );
  XOR U3802 ( .A(n3939), .B(n3931), .Z(n3923) );
  XOR U3803 ( .A(n3720), .B(n3940), .Z(n3931) );
  IV U3804 ( .A(n3719), .Z(n3940) );
  XNOR U3805 ( .A(n3716), .B(n3941), .Z(n3719) );
  XOR U3806 ( .A(n3942), .B(n3943), .Z(n3716) );
  ANDN U3807 ( .A(n3944), .B(n3945), .Z(n3943) );
  XNOR U3808 ( .A(n3942), .B(n3946), .Z(n3944) );
  XOR U3809 ( .A(n3727), .B(n3947), .Z(n3720) );
  IV U3810 ( .A(n3726), .Z(n3947) );
  XNOR U3811 ( .A(n3723), .B(n3948), .Z(n3726) );
  XOR U3812 ( .A(n3949), .B(n3950), .Z(n3723) );
  ANDN U3813 ( .A(n3951), .B(n3952), .Z(n3950) );
  XNOR U3814 ( .A(n3949), .B(n3953), .Z(n3951) );
  XOR U3815 ( .A(n3734), .B(n3954), .Z(n3727) );
  IV U3816 ( .A(n3733), .Z(n3954) );
  XNOR U3817 ( .A(n3730), .B(n3955), .Z(n3733) );
  XOR U3818 ( .A(n3956), .B(n3957), .Z(n3730) );
  ANDN U3819 ( .A(n3958), .B(n3959), .Z(n3957) );
  XNOR U3820 ( .A(n3956), .B(n3960), .Z(n3958) );
  XOR U3821 ( .A(n3741), .B(n3961), .Z(n3734) );
  IV U3822 ( .A(n3740), .Z(n3961) );
  XNOR U3823 ( .A(n3737), .B(n3962), .Z(n3740) );
  XOR U3824 ( .A(n3963), .B(n3964), .Z(n3737) );
  ANDN U3825 ( .A(n3965), .B(n3966), .Z(n3964) );
  XNOR U3826 ( .A(n3963), .B(n3967), .Z(n3965) );
  XOR U3827 ( .A(n3748), .B(n3968), .Z(n3741) );
  IV U3828 ( .A(n3747), .Z(n3968) );
  XNOR U3829 ( .A(n3744), .B(n3969), .Z(n3747) );
  XOR U3830 ( .A(n3970), .B(n3971), .Z(n3744) );
  ANDN U3831 ( .A(n3972), .B(n3973), .Z(n3971) );
  XNOR U3832 ( .A(n3970), .B(n3974), .Z(n3972) );
  XOR U3833 ( .A(n3755), .B(n3975), .Z(n3748) );
  IV U3834 ( .A(n3754), .Z(n3975) );
  XNOR U3835 ( .A(n3751), .B(n3976), .Z(n3754) );
  XOR U3836 ( .A(n3977), .B(n3978), .Z(n3751) );
  ANDN U3837 ( .A(n3979), .B(n3980), .Z(n3978) );
  XNOR U3838 ( .A(n3977), .B(n3981), .Z(n3979) );
  XOR U3839 ( .A(n3762), .B(n3982), .Z(n3755) );
  IV U3840 ( .A(n3761), .Z(n3982) );
  XNOR U3841 ( .A(n3758), .B(n3983), .Z(n3761) );
  XOR U3842 ( .A(n3984), .B(n3985), .Z(n3758) );
  ANDN U3843 ( .A(n3986), .B(n3987), .Z(n3985) );
  XNOR U3844 ( .A(n3984), .B(n3988), .Z(n3986) );
  XOR U3845 ( .A(n3769), .B(n3989), .Z(n3762) );
  IV U3846 ( .A(n3768), .Z(n3989) );
  XNOR U3847 ( .A(n3765), .B(n3990), .Z(n3768) );
  XOR U3848 ( .A(n3991), .B(n3992), .Z(n3765) );
  ANDN U3849 ( .A(n3993), .B(n3994), .Z(n3992) );
  XNOR U3850 ( .A(n3991), .B(n3995), .Z(n3993) );
  XOR U3851 ( .A(n3776), .B(n3996), .Z(n3769) );
  IV U3852 ( .A(n3775), .Z(n3996) );
  XNOR U3853 ( .A(n3772), .B(n3997), .Z(n3775) );
  XOR U3854 ( .A(n3998), .B(n3999), .Z(n3772) );
  ANDN U3855 ( .A(n4000), .B(n4001), .Z(n3999) );
  XNOR U3856 ( .A(n3998), .B(n4002), .Z(n4000) );
  XOR U3857 ( .A(n3783), .B(n4003), .Z(n3776) );
  IV U3858 ( .A(n3782), .Z(n4003) );
  XNOR U3859 ( .A(n3779), .B(n4004), .Z(n3782) );
  XOR U3860 ( .A(n4005), .B(n4006), .Z(n3779) );
  ANDN U3861 ( .A(n4007), .B(n4008), .Z(n4006) );
  XNOR U3862 ( .A(n4005), .B(n4009), .Z(n4007) );
  XOR U3863 ( .A(n3790), .B(n4010), .Z(n3783) );
  IV U3864 ( .A(n3789), .Z(n4010) );
  XNOR U3865 ( .A(n3786), .B(n4011), .Z(n3789) );
  XOR U3866 ( .A(n4012), .B(n4013), .Z(n3786) );
  ANDN U3867 ( .A(n4014), .B(n4015), .Z(n4013) );
  XNOR U3868 ( .A(n4012), .B(n4016), .Z(n4014) );
  XOR U3869 ( .A(n3797), .B(n4017), .Z(n3790) );
  IV U3870 ( .A(n3796), .Z(n4017) );
  XNOR U3871 ( .A(n3793), .B(n4018), .Z(n3796) );
  XOR U3872 ( .A(n4019), .B(n4020), .Z(n3793) );
  ANDN U3873 ( .A(n4021), .B(n4022), .Z(n4020) );
  XNOR U3874 ( .A(n4019), .B(n4023), .Z(n4021) );
  XOR U3875 ( .A(n3804), .B(n4024), .Z(n3797) );
  IV U3876 ( .A(n3803), .Z(n4024) );
  XNOR U3877 ( .A(n3800), .B(n4025), .Z(n3803) );
  XOR U3878 ( .A(n4026), .B(n4027), .Z(n3800) );
  ANDN U3879 ( .A(n4028), .B(n4029), .Z(n4027) );
  XNOR U3880 ( .A(n4026), .B(n4030), .Z(n4028) );
  XOR U3881 ( .A(n3811), .B(n4031), .Z(n3804) );
  IV U3882 ( .A(n3810), .Z(n4031) );
  XNOR U3883 ( .A(n3807), .B(n4032), .Z(n3810) );
  XOR U3884 ( .A(n4033), .B(n4034), .Z(n3807) );
  ANDN U3885 ( .A(n4035), .B(n4036), .Z(n4034) );
  XNOR U3886 ( .A(n4033), .B(n4037), .Z(n4035) );
  XOR U3887 ( .A(n3818), .B(n4038), .Z(n3811) );
  IV U3888 ( .A(n3817), .Z(n4038) );
  XNOR U3889 ( .A(n3814), .B(n4039), .Z(n3817) );
  XOR U3890 ( .A(n4040), .B(n4041), .Z(n3814) );
  ANDN U3891 ( .A(n4042), .B(n4043), .Z(n4041) );
  XNOR U3892 ( .A(n4040), .B(n4044), .Z(n4042) );
  XOR U3893 ( .A(n3824), .B(n4045), .Z(n3818) );
  IV U3894 ( .A(n3823), .Z(n4045) );
  XNOR U3895 ( .A(n3820), .B(n4046), .Z(n3823) );
  XOR U3896 ( .A(n4047), .B(n4048), .Z(n3820) );
  ANDN U3897 ( .A(n4049), .B(n4050), .Z(n4048) );
  XNOR U3898 ( .A(n4047), .B(n4051), .Z(n4049) );
  XOR U3899 ( .A(n3830), .B(n4052), .Z(n3824) );
  IV U3900 ( .A(n3829), .Z(n4052) );
  XNOR U3901 ( .A(n3826), .B(n4039), .Z(n3829) );
  AND U3902 ( .A(n4525), .B(n3593), .Z(n4039) );
  XOR U3903 ( .A(n4053), .B(n4054), .Z(n3826) );
  ANDN U3904 ( .A(n4055), .B(n4056), .Z(n4054) );
  XNOR U3905 ( .A(n4053), .B(n4057), .Z(n4055) );
  XOR U3906 ( .A(n3836), .B(n4058), .Z(n3830) );
  IV U3907 ( .A(n3835), .Z(n4058) );
  XNOR U3908 ( .A(n3832), .B(n4032), .Z(n3835) );
  AND U3909 ( .A(n5030), .B(n3166), .Z(n4032) );
  XOR U3910 ( .A(n4059), .B(n4060), .Z(n3832) );
  ANDN U3911 ( .A(n4061), .B(n4062), .Z(n4060) );
  XNOR U3912 ( .A(n4059), .B(n4063), .Z(n4061) );
  XOR U3913 ( .A(n3842), .B(n4064), .Z(n3836) );
  IV U3914 ( .A(n3841), .Z(n4064) );
  XNOR U3915 ( .A(n3838), .B(n4025), .Z(n3841) );
  AND U3916 ( .A(n5561), .B(n2765), .Z(n4025) );
  XOR U3917 ( .A(n4065), .B(n4066), .Z(n3838) );
  ANDN U3918 ( .A(n4067), .B(n4068), .Z(n4066) );
  XNOR U3919 ( .A(n4065), .B(n4069), .Z(n4067) );
  XOR U3920 ( .A(n3848), .B(n4070), .Z(n3842) );
  IV U3921 ( .A(n3847), .Z(n4070) );
  XNOR U3922 ( .A(n3844), .B(n4018), .Z(n3847) );
  AND U3923 ( .A(n6118), .B(n2396), .Z(n4018) );
  XOR U3924 ( .A(n4071), .B(n4072), .Z(n3844) );
  ANDN U3925 ( .A(n4073), .B(n4074), .Z(n4072) );
  XNOR U3926 ( .A(n4071), .B(n4075), .Z(n4073) );
  XOR U3927 ( .A(n3854), .B(n4076), .Z(n3848) );
  IV U3928 ( .A(n3853), .Z(n4076) );
  XNOR U3929 ( .A(n3850), .B(n4011), .Z(n3853) );
  AND U3930 ( .A(n6688), .B(n2053), .Z(n4011) );
  XOR U3931 ( .A(n4077), .B(n4078), .Z(n3850) );
  ANDN U3932 ( .A(n4079), .B(n4080), .Z(n4078) );
  XNOR U3933 ( .A(n4077), .B(n4081), .Z(n4079) );
  XOR U3934 ( .A(n3860), .B(n4082), .Z(n3854) );
  IV U3935 ( .A(n3859), .Z(n4082) );
  XNOR U3936 ( .A(n3856), .B(n4004), .Z(n3859) );
  AND U3937 ( .A(n7241), .B(n1737), .Z(n4004) );
  XOR U3938 ( .A(n4083), .B(n4084), .Z(n3856) );
  ANDN U3939 ( .A(n4085), .B(n4086), .Z(n4084) );
  XNOR U3940 ( .A(n4083), .B(n4087), .Z(n4085) );
  XOR U3941 ( .A(n3866), .B(n4088), .Z(n3860) );
  IV U3942 ( .A(n3865), .Z(n4088) );
  XNOR U3943 ( .A(n3862), .B(n3997), .Z(n3865) );
  AND U3944 ( .A(n7770), .B(n1448), .Z(n3997) );
  XOR U3945 ( .A(n4089), .B(n4090), .Z(n3862) );
  ANDN U3946 ( .A(n4091), .B(n4092), .Z(n4090) );
  XNOR U3947 ( .A(n4089), .B(n4093), .Z(n4091) );
  XOR U3948 ( .A(n3872), .B(n4094), .Z(n3866) );
  IV U3949 ( .A(n3871), .Z(n4094) );
  XNOR U3950 ( .A(n3868), .B(n3990), .Z(n3871) );
  AND U3951 ( .A(n8272), .B(n1185), .Z(n3990) );
  XOR U3952 ( .A(n4095), .B(n4096), .Z(n3868) );
  ANDN U3953 ( .A(n4097), .B(n4098), .Z(n4096) );
  XNOR U3954 ( .A(n4095), .B(n4099), .Z(n4097) );
  XOR U3955 ( .A(n3878), .B(n4100), .Z(n3872) );
  IV U3956 ( .A(n3877), .Z(n4100) );
  XNOR U3957 ( .A(n3874), .B(n3983), .Z(n3877) );
  AND U3958 ( .A(n8748), .B(n948), .Z(n3983) );
  XOR U3959 ( .A(n4101), .B(n4102), .Z(n3874) );
  ANDN U3960 ( .A(n4103), .B(n4104), .Z(n4102) );
  XNOR U3961 ( .A(n4101), .B(n4105), .Z(n4103) );
  XOR U3962 ( .A(n3884), .B(n4106), .Z(n3878) );
  IV U3963 ( .A(n3883), .Z(n4106) );
  XNOR U3964 ( .A(n3880), .B(n3976), .Z(n3883) );
  AND U3965 ( .A(n9198), .B(n736), .Z(n3976) );
  XOR U3966 ( .A(n4107), .B(n4108), .Z(n3880) );
  ANDN U3967 ( .A(n4109), .B(n4110), .Z(n4108) );
  XNOR U3968 ( .A(n4107), .B(n4111), .Z(n4109) );
  XOR U3969 ( .A(n3890), .B(n4112), .Z(n3884) );
  IV U3970 ( .A(n3889), .Z(n4112) );
  XNOR U3971 ( .A(n3886), .B(n3969), .Z(n3889) );
  AND U3972 ( .A(n9621), .B(n552), .Z(n3969) );
  XOR U3973 ( .A(n4113), .B(n4114), .Z(n3886) );
  ANDN U3974 ( .A(n4115), .B(n4116), .Z(n4114) );
  XNOR U3975 ( .A(n4113), .B(n4117), .Z(n4115) );
  XOR U3976 ( .A(n3896), .B(n4118), .Z(n3890) );
  IV U3977 ( .A(n3895), .Z(n4118) );
  XNOR U3978 ( .A(n3892), .B(n3962), .Z(n3895) );
  AND U3979 ( .A(n10017), .B(n395), .Z(n3962) );
  XOR U3980 ( .A(n4119), .B(n4120), .Z(n3892) );
  ANDN U3981 ( .A(n4121), .B(n4122), .Z(n4120) );
  XNOR U3982 ( .A(n4119), .B(n4123), .Z(n4121) );
  XOR U3983 ( .A(n3902), .B(n4124), .Z(n3896) );
  IV U3984 ( .A(n3901), .Z(n4124) );
  XNOR U3985 ( .A(n3898), .B(n3955), .Z(n3901) );
  AND U3986 ( .A(n10387), .B(n264), .Z(n3955) );
  XOR U3987 ( .A(n4125), .B(n4126), .Z(n3898) );
  ANDN U3988 ( .A(n4127), .B(n4128), .Z(n4126) );
  XNOR U3989 ( .A(n4125), .B(n4129), .Z(n4127) );
  XOR U3990 ( .A(n3908), .B(n4130), .Z(n3902) );
  IV U3991 ( .A(n3907), .Z(n4130) );
  XNOR U3992 ( .A(n3904), .B(n3948), .Z(n3907) );
  AND U3993 ( .A(n10731), .B(n159), .Z(n3948) );
  XOR U3994 ( .A(n4131), .B(n4132), .Z(n3904) );
  ANDN U3995 ( .A(n4133), .B(n4134), .Z(n4132) );
  XNOR U3996 ( .A(n4131), .B(n4135), .Z(n4133) );
  XOR U3997 ( .A(n3915), .B(n4136), .Z(n3908) );
  IV U3998 ( .A(n3914), .Z(n4136) );
  XNOR U3999 ( .A(n3911), .B(n3941), .Z(n3914) );
  AND U4000 ( .A(n11049), .B(n80), .Z(n3941) );
  XOR U4001 ( .A(n4137), .B(n4138), .Z(n3911) );
  ANDN U4002 ( .A(n4139), .B(n4140), .Z(n4138) );
  XNOR U4003 ( .A(n4137), .B(n4141), .Z(n4139) );
  XOR U4004 ( .A(n3920), .B(n4142), .Z(n3915) );
  IV U4005 ( .A(n3919), .Z(n4142) );
  XNOR U4006 ( .A(n3916), .B(n4143), .Z(n3919) );
  AND U4007 ( .A(n42), .B(n11341), .Z(n4143) );
  XOR U4008 ( .A(n4144), .B(n4145), .Z(n3916) );
  ANDN U4009 ( .A(n4146), .B(n4147), .Z(n4145) );
  XNOR U4010 ( .A(n4144), .B(n4148), .Z(n4146) );
  XNOR U4011 ( .A(n4149), .B(n4150), .Z(n3920) );
  ANDN U4012 ( .A(n4151), .B(n4152), .Z(n4150) );
  XNOR U4013 ( .A(n4149), .B(n4153), .Z(n4151) );
  XNOR U4014 ( .A(n3929), .B(n3921), .Z(n3939) );
  XOR U4015 ( .A(n4154), .B(n4155), .Z(n3921) );
  AND U4016 ( .A(n4156), .B(n4157), .Z(n4155) );
  XNOR U4017 ( .A(n4158), .B(n4154), .Z(n4157) );
  XOR U4018 ( .A(n3927), .B(n4159), .Z(n3929) );
  ANDN U4019 ( .A(n11341), .B(n43), .Z(n4159) );
  XOR U4020 ( .A(n4160), .B(n4161), .Z(n3927) );
  AND U4021 ( .A(n4162), .B(n4163), .Z(n4161) );
  XNOR U4022 ( .A(n4160), .B(n4164), .Z(n4163) );
  XOR U4023 ( .A(n3925), .B(n3935), .Z(n3938) );
  XOR U4024 ( .A(n4165), .B(n4166), .Z(n3925) );
  IV U4025 ( .A(n4167), .Z(n4166) );
  XOR U4026 ( .A(n4168), .B(n4169), .Z(n3935) );
  AND U4027 ( .A(n4168), .B(n4170), .Z(n4169) );
  XOR U4028 ( .A(n4171), .B(n4156), .Z(n4170) );
  XOR U4029 ( .A(n4172), .B(n4164), .Z(n4156) );
  XOR U4030 ( .A(n3946), .B(n4173), .Z(n4164) );
  IV U4031 ( .A(n3945), .Z(n4173) );
  XNOR U4032 ( .A(n3942), .B(n4174), .Z(n3945) );
  XOR U4033 ( .A(n4175), .B(n4176), .Z(n3942) );
  ANDN U4034 ( .A(n4177), .B(n4178), .Z(n4176) );
  XNOR U4035 ( .A(n4175), .B(n4179), .Z(n4177) );
  XOR U4036 ( .A(n3953), .B(n4180), .Z(n3946) );
  IV U4037 ( .A(n3952), .Z(n4180) );
  XNOR U4038 ( .A(n3949), .B(n4181), .Z(n3952) );
  XOR U4039 ( .A(n4182), .B(n4183), .Z(n3949) );
  ANDN U4040 ( .A(n4184), .B(n4185), .Z(n4183) );
  XNOR U4041 ( .A(n4182), .B(n4186), .Z(n4184) );
  XOR U4042 ( .A(n3960), .B(n4187), .Z(n3953) );
  IV U4043 ( .A(n3959), .Z(n4187) );
  XNOR U4044 ( .A(n3956), .B(n4188), .Z(n3959) );
  XOR U4045 ( .A(n4189), .B(n4190), .Z(n3956) );
  ANDN U4046 ( .A(n4191), .B(n4192), .Z(n4190) );
  XNOR U4047 ( .A(n4189), .B(n4193), .Z(n4191) );
  XOR U4048 ( .A(n3967), .B(n4194), .Z(n3960) );
  IV U4049 ( .A(n3966), .Z(n4194) );
  XNOR U4050 ( .A(n3963), .B(n4195), .Z(n3966) );
  XOR U4051 ( .A(n4196), .B(n4197), .Z(n3963) );
  ANDN U4052 ( .A(n4198), .B(n4199), .Z(n4197) );
  XNOR U4053 ( .A(n4196), .B(n4200), .Z(n4198) );
  XOR U4054 ( .A(n3974), .B(n4201), .Z(n3967) );
  IV U4055 ( .A(n3973), .Z(n4201) );
  XNOR U4056 ( .A(n3970), .B(n4202), .Z(n3973) );
  XOR U4057 ( .A(n4203), .B(n4204), .Z(n3970) );
  ANDN U4058 ( .A(n4205), .B(n4206), .Z(n4204) );
  XNOR U4059 ( .A(n4203), .B(n4207), .Z(n4205) );
  XOR U4060 ( .A(n3981), .B(n4208), .Z(n3974) );
  IV U4061 ( .A(n3980), .Z(n4208) );
  XNOR U4062 ( .A(n3977), .B(n4209), .Z(n3980) );
  XOR U4063 ( .A(n4210), .B(n4211), .Z(n3977) );
  ANDN U4064 ( .A(n4212), .B(n4213), .Z(n4211) );
  XNOR U4065 ( .A(n4210), .B(n4214), .Z(n4212) );
  XOR U4066 ( .A(n3988), .B(n4215), .Z(n3981) );
  IV U4067 ( .A(n3987), .Z(n4215) );
  XNOR U4068 ( .A(n3984), .B(n4216), .Z(n3987) );
  XOR U4069 ( .A(n4217), .B(n4218), .Z(n3984) );
  ANDN U4070 ( .A(n4219), .B(n4220), .Z(n4218) );
  XNOR U4071 ( .A(n4217), .B(n4221), .Z(n4219) );
  XOR U4072 ( .A(n3995), .B(n4222), .Z(n3988) );
  IV U4073 ( .A(n3994), .Z(n4222) );
  XNOR U4074 ( .A(n3991), .B(n4223), .Z(n3994) );
  XOR U4075 ( .A(n4224), .B(n4225), .Z(n3991) );
  ANDN U4076 ( .A(n4226), .B(n4227), .Z(n4225) );
  XNOR U4077 ( .A(n4224), .B(n4228), .Z(n4226) );
  XOR U4078 ( .A(n4002), .B(n4229), .Z(n3995) );
  IV U4079 ( .A(n4001), .Z(n4229) );
  XNOR U4080 ( .A(n3998), .B(n4230), .Z(n4001) );
  XOR U4081 ( .A(n4231), .B(n4232), .Z(n3998) );
  ANDN U4082 ( .A(n4233), .B(n4234), .Z(n4232) );
  XNOR U4083 ( .A(n4231), .B(n4235), .Z(n4233) );
  XOR U4084 ( .A(n4009), .B(n4236), .Z(n4002) );
  IV U4085 ( .A(n4008), .Z(n4236) );
  XNOR U4086 ( .A(n4005), .B(n4237), .Z(n4008) );
  XOR U4087 ( .A(n4238), .B(n4239), .Z(n4005) );
  ANDN U4088 ( .A(n4240), .B(n4241), .Z(n4239) );
  XNOR U4089 ( .A(n4238), .B(n4242), .Z(n4240) );
  XOR U4090 ( .A(n4016), .B(n4243), .Z(n4009) );
  IV U4091 ( .A(n4015), .Z(n4243) );
  XNOR U4092 ( .A(n4012), .B(n4244), .Z(n4015) );
  XOR U4093 ( .A(n4245), .B(n4246), .Z(n4012) );
  ANDN U4094 ( .A(n4247), .B(n4248), .Z(n4246) );
  XNOR U4095 ( .A(n4245), .B(n4249), .Z(n4247) );
  XOR U4096 ( .A(n4023), .B(n4250), .Z(n4016) );
  IV U4097 ( .A(n4022), .Z(n4250) );
  XNOR U4098 ( .A(n4019), .B(n4251), .Z(n4022) );
  XOR U4099 ( .A(n4252), .B(n4253), .Z(n4019) );
  ANDN U4100 ( .A(n4254), .B(n4255), .Z(n4253) );
  XNOR U4101 ( .A(n4252), .B(n4256), .Z(n4254) );
  XOR U4102 ( .A(n4030), .B(n4257), .Z(n4023) );
  IV U4103 ( .A(n4029), .Z(n4257) );
  XNOR U4104 ( .A(n4026), .B(n4258), .Z(n4029) );
  XOR U4105 ( .A(n4259), .B(n4260), .Z(n4026) );
  ANDN U4106 ( .A(n4261), .B(n4262), .Z(n4260) );
  XNOR U4107 ( .A(n4259), .B(n4263), .Z(n4261) );
  XOR U4108 ( .A(n4037), .B(n4264), .Z(n4030) );
  IV U4109 ( .A(n4036), .Z(n4264) );
  XNOR U4110 ( .A(n4033), .B(n4265), .Z(n4036) );
  XOR U4111 ( .A(n4266), .B(n4267), .Z(n4033) );
  ANDN U4112 ( .A(n4268), .B(n4269), .Z(n4267) );
  XNOR U4113 ( .A(n4266), .B(n4270), .Z(n4268) );
  XOR U4114 ( .A(n4044), .B(n4271), .Z(n4037) );
  IV U4115 ( .A(n4043), .Z(n4271) );
  XNOR U4116 ( .A(n4040), .B(n4272), .Z(n4043) );
  XOR U4117 ( .A(n4273), .B(n4274), .Z(n4040) );
  ANDN U4118 ( .A(n4275), .B(n4276), .Z(n4274) );
  XNOR U4119 ( .A(n4273), .B(n4277), .Z(n4275) );
  XOR U4120 ( .A(n4051), .B(n4278), .Z(n4044) );
  IV U4121 ( .A(n4050), .Z(n4278) );
  XNOR U4122 ( .A(n4047), .B(n4279), .Z(n4050) );
  XOR U4123 ( .A(n4280), .B(n4281), .Z(n4047) );
  ANDN U4124 ( .A(n4282), .B(n4283), .Z(n4281) );
  XNOR U4125 ( .A(n4280), .B(n4284), .Z(n4282) );
  XOR U4126 ( .A(n4057), .B(n4285), .Z(n4051) );
  IV U4127 ( .A(n4056), .Z(n4285) );
  XNOR U4128 ( .A(n4053), .B(n4279), .Z(n4056) );
  AND U4129 ( .A(n4525), .B(n4046), .Z(n4279) );
  XOR U4130 ( .A(n4286), .B(n4287), .Z(n4053) );
  ANDN U4131 ( .A(n4288), .B(n4289), .Z(n4287) );
  XNOR U4132 ( .A(n4286), .B(n4290), .Z(n4288) );
  XOR U4133 ( .A(n4063), .B(n4291), .Z(n4057) );
  IV U4134 ( .A(n4062), .Z(n4291) );
  XNOR U4135 ( .A(n4059), .B(n4272), .Z(n4062) );
  AND U4136 ( .A(n5030), .B(n3593), .Z(n4272) );
  XOR U4137 ( .A(n4292), .B(n4293), .Z(n4059) );
  ANDN U4138 ( .A(n4294), .B(n4295), .Z(n4293) );
  XNOR U4139 ( .A(n4292), .B(n4296), .Z(n4294) );
  XOR U4140 ( .A(n4069), .B(n4297), .Z(n4063) );
  IV U4141 ( .A(n4068), .Z(n4297) );
  XNOR U4142 ( .A(n4065), .B(n4265), .Z(n4068) );
  AND U4143 ( .A(n5561), .B(n3166), .Z(n4265) );
  XOR U4144 ( .A(n4298), .B(n4299), .Z(n4065) );
  ANDN U4145 ( .A(n4300), .B(n4301), .Z(n4299) );
  XNOR U4146 ( .A(n4298), .B(n4302), .Z(n4300) );
  XOR U4147 ( .A(n4075), .B(n4303), .Z(n4069) );
  IV U4148 ( .A(n4074), .Z(n4303) );
  XNOR U4149 ( .A(n4071), .B(n4258), .Z(n4074) );
  AND U4150 ( .A(n6118), .B(n2765), .Z(n4258) );
  XOR U4151 ( .A(n4304), .B(n4305), .Z(n4071) );
  ANDN U4152 ( .A(n4306), .B(n4307), .Z(n4305) );
  XNOR U4153 ( .A(n4304), .B(n4308), .Z(n4306) );
  XOR U4154 ( .A(n4081), .B(n4309), .Z(n4075) );
  IV U4155 ( .A(n4080), .Z(n4309) );
  XNOR U4156 ( .A(n4077), .B(n4251), .Z(n4080) );
  AND U4157 ( .A(n6688), .B(n2396), .Z(n4251) );
  XOR U4158 ( .A(n4310), .B(n4311), .Z(n4077) );
  ANDN U4159 ( .A(n4312), .B(n4313), .Z(n4311) );
  XNOR U4160 ( .A(n4310), .B(n4314), .Z(n4312) );
  XOR U4161 ( .A(n4087), .B(n4315), .Z(n4081) );
  IV U4162 ( .A(n4086), .Z(n4315) );
  XNOR U4163 ( .A(n4083), .B(n4244), .Z(n4086) );
  AND U4164 ( .A(n7241), .B(n2053), .Z(n4244) );
  XOR U4165 ( .A(n4316), .B(n4317), .Z(n4083) );
  ANDN U4166 ( .A(n4318), .B(n4319), .Z(n4317) );
  XNOR U4167 ( .A(n4316), .B(n4320), .Z(n4318) );
  XOR U4168 ( .A(n4093), .B(n4321), .Z(n4087) );
  IV U4169 ( .A(n4092), .Z(n4321) );
  XNOR U4170 ( .A(n4089), .B(n4237), .Z(n4092) );
  AND U4171 ( .A(n7770), .B(n1737), .Z(n4237) );
  XOR U4172 ( .A(n4322), .B(n4323), .Z(n4089) );
  ANDN U4173 ( .A(n4324), .B(n4325), .Z(n4323) );
  XNOR U4174 ( .A(n4322), .B(n4326), .Z(n4324) );
  XOR U4175 ( .A(n4099), .B(n4327), .Z(n4093) );
  IV U4176 ( .A(n4098), .Z(n4327) );
  XNOR U4177 ( .A(n4095), .B(n4230), .Z(n4098) );
  AND U4178 ( .A(n8272), .B(n1448), .Z(n4230) );
  XOR U4179 ( .A(n4328), .B(n4329), .Z(n4095) );
  ANDN U4180 ( .A(n4330), .B(n4331), .Z(n4329) );
  XNOR U4181 ( .A(n4328), .B(n4332), .Z(n4330) );
  XOR U4182 ( .A(n4105), .B(n4333), .Z(n4099) );
  IV U4183 ( .A(n4104), .Z(n4333) );
  XNOR U4184 ( .A(n4101), .B(n4223), .Z(n4104) );
  AND U4185 ( .A(n8748), .B(n1185), .Z(n4223) );
  XOR U4186 ( .A(n4334), .B(n4335), .Z(n4101) );
  ANDN U4187 ( .A(n4336), .B(n4337), .Z(n4335) );
  XNOR U4188 ( .A(n4334), .B(n4338), .Z(n4336) );
  XOR U4189 ( .A(n4111), .B(n4339), .Z(n4105) );
  IV U4190 ( .A(n4110), .Z(n4339) );
  XNOR U4191 ( .A(n4107), .B(n4216), .Z(n4110) );
  AND U4192 ( .A(n9198), .B(n948), .Z(n4216) );
  XOR U4193 ( .A(n4340), .B(n4341), .Z(n4107) );
  ANDN U4194 ( .A(n4342), .B(n4343), .Z(n4341) );
  XNOR U4195 ( .A(n4340), .B(n4344), .Z(n4342) );
  XOR U4196 ( .A(n4117), .B(n4345), .Z(n4111) );
  IV U4197 ( .A(n4116), .Z(n4345) );
  XNOR U4198 ( .A(n4113), .B(n4209), .Z(n4116) );
  AND U4199 ( .A(n9621), .B(n736), .Z(n4209) );
  XOR U4200 ( .A(n4346), .B(n4347), .Z(n4113) );
  ANDN U4201 ( .A(n4348), .B(n4349), .Z(n4347) );
  XNOR U4202 ( .A(n4346), .B(n4350), .Z(n4348) );
  XOR U4203 ( .A(n4123), .B(n4351), .Z(n4117) );
  IV U4204 ( .A(n4122), .Z(n4351) );
  XNOR U4205 ( .A(n4119), .B(n4202), .Z(n4122) );
  AND U4206 ( .A(n10017), .B(n552), .Z(n4202) );
  XOR U4207 ( .A(n4352), .B(n4353), .Z(n4119) );
  ANDN U4208 ( .A(n4354), .B(n4355), .Z(n4353) );
  XNOR U4209 ( .A(n4352), .B(n4356), .Z(n4354) );
  XOR U4210 ( .A(n4129), .B(n4357), .Z(n4123) );
  IV U4211 ( .A(n4128), .Z(n4357) );
  XNOR U4212 ( .A(n4125), .B(n4195), .Z(n4128) );
  AND U4213 ( .A(n10387), .B(n395), .Z(n4195) );
  XOR U4214 ( .A(n4358), .B(n4359), .Z(n4125) );
  ANDN U4215 ( .A(n4360), .B(n4361), .Z(n4359) );
  XNOR U4216 ( .A(n4358), .B(n4362), .Z(n4360) );
  XOR U4217 ( .A(n4135), .B(n4363), .Z(n4129) );
  IV U4218 ( .A(n4134), .Z(n4363) );
  XNOR U4219 ( .A(n4131), .B(n4188), .Z(n4134) );
  AND U4220 ( .A(n10731), .B(n264), .Z(n4188) );
  XOR U4221 ( .A(n4364), .B(n4365), .Z(n4131) );
  ANDN U4222 ( .A(n4366), .B(n4367), .Z(n4365) );
  XNOR U4223 ( .A(n4364), .B(n4368), .Z(n4366) );
  XOR U4224 ( .A(n4141), .B(n4369), .Z(n4135) );
  IV U4225 ( .A(n4140), .Z(n4369) );
  XNOR U4226 ( .A(n4137), .B(n4181), .Z(n4140) );
  AND U4227 ( .A(n11049), .B(n159), .Z(n4181) );
  XOR U4228 ( .A(n4370), .B(n4371), .Z(n4137) );
  ANDN U4229 ( .A(n4372), .B(n4373), .Z(n4371) );
  XNOR U4230 ( .A(n4370), .B(n4374), .Z(n4372) );
  XOR U4231 ( .A(n4148), .B(n4375), .Z(n4141) );
  IV U4232 ( .A(n4147), .Z(n4375) );
  XNOR U4233 ( .A(n4144), .B(n4174), .Z(n4147) );
  AND U4234 ( .A(n11341), .B(n80), .Z(n4174) );
  XOR U4235 ( .A(n4376), .B(n4377), .Z(n4144) );
  ANDN U4236 ( .A(n4378), .B(n4379), .Z(n4377) );
  XNOR U4237 ( .A(n4376), .B(n4380), .Z(n4378) );
  XOR U4238 ( .A(n4153), .B(n4381), .Z(n4148) );
  IV U4239 ( .A(n4152), .Z(n4381) );
  XNOR U4240 ( .A(n4149), .B(n4382), .Z(n4152) );
  AND U4241 ( .A(n42), .B(n11607), .Z(n4382) );
  XOR U4242 ( .A(n4383), .B(n4384), .Z(n4149) );
  ANDN U4243 ( .A(n4385), .B(n4386), .Z(n4384) );
  XNOR U4244 ( .A(n4383), .B(n4387), .Z(n4385) );
  XNOR U4245 ( .A(n4388), .B(n4389), .Z(n4153) );
  ANDN U4246 ( .A(n4390), .B(n4391), .Z(n4389) );
  XNOR U4247 ( .A(n4388), .B(n4392), .Z(n4390) );
  XNOR U4248 ( .A(n4162), .B(n4154), .Z(n4172) );
  XOR U4249 ( .A(n4393), .B(n4394), .Z(n4154) );
  AND U4250 ( .A(n4395), .B(n4396), .Z(n4394) );
  XNOR U4251 ( .A(n4397), .B(n4393), .Z(n4396) );
  XOR U4252 ( .A(n4160), .B(n4398), .Z(n4162) );
  ANDN U4253 ( .A(n11607), .B(n43), .Z(n4398) );
  XOR U4254 ( .A(n4399), .B(n4400), .Z(n4160) );
  AND U4255 ( .A(n4401), .B(n4402), .Z(n4400) );
  XNOR U4256 ( .A(n4399), .B(n4403), .Z(n4402) );
  XOR U4257 ( .A(n4158), .B(n4168), .Z(n4171) );
  XOR U4258 ( .A(n4404), .B(n4405), .Z(n4158) );
  IV U4259 ( .A(n4406), .Z(n4405) );
  XOR U4260 ( .A(n4407), .B(n4408), .Z(n4168) );
  AND U4261 ( .A(n4407), .B(n4409), .Z(n4408) );
  XOR U4262 ( .A(n4410), .B(n4395), .Z(n4409) );
  XOR U4263 ( .A(n4411), .B(n4403), .Z(n4395) );
  XOR U4264 ( .A(n4179), .B(n4412), .Z(n4403) );
  IV U4265 ( .A(n4178), .Z(n4412) );
  XNOR U4266 ( .A(n4175), .B(n4413), .Z(n4178) );
  XOR U4267 ( .A(n4414), .B(n4415), .Z(n4175) );
  ANDN U4268 ( .A(n4416), .B(n4417), .Z(n4415) );
  XNOR U4269 ( .A(n4414), .B(n4418), .Z(n4416) );
  XOR U4270 ( .A(n4186), .B(n4419), .Z(n4179) );
  IV U4271 ( .A(n4185), .Z(n4419) );
  XNOR U4272 ( .A(n4182), .B(n4420), .Z(n4185) );
  XOR U4273 ( .A(n4421), .B(n4422), .Z(n4182) );
  ANDN U4274 ( .A(n4423), .B(n4424), .Z(n4422) );
  XNOR U4275 ( .A(n4421), .B(n4425), .Z(n4423) );
  XOR U4276 ( .A(n4193), .B(n4426), .Z(n4186) );
  IV U4277 ( .A(n4192), .Z(n4426) );
  XNOR U4278 ( .A(n4189), .B(n4427), .Z(n4192) );
  XOR U4279 ( .A(n4428), .B(n4429), .Z(n4189) );
  ANDN U4280 ( .A(n4430), .B(n4431), .Z(n4429) );
  XNOR U4281 ( .A(n4428), .B(n4432), .Z(n4430) );
  XOR U4282 ( .A(n4200), .B(n4433), .Z(n4193) );
  IV U4283 ( .A(n4199), .Z(n4433) );
  XNOR U4284 ( .A(n4196), .B(n4434), .Z(n4199) );
  XOR U4285 ( .A(n4435), .B(n4436), .Z(n4196) );
  ANDN U4286 ( .A(n4437), .B(n4438), .Z(n4436) );
  XNOR U4287 ( .A(n4435), .B(n4439), .Z(n4437) );
  XOR U4288 ( .A(n4207), .B(n4440), .Z(n4200) );
  IV U4289 ( .A(n4206), .Z(n4440) );
  XNOR U4290 ( .A(n4203), .B(n4441), .Z(n4206) );
  XOR U4291 ( .A(n4442), .B(n4443), .Z(n4203) );
  ANDN U4292 ( .A(n4444), .B(n4445), .Z(n4443) );
  XNOR U4293 ( .A(n4442), .B(n4446), .Z(n4444) );
  XOR U4294 ( .A(n4214), .B(n4447), .Z(n4207) );
  IV U4295 ( .A(n4213), .Z(n4447) );
  XNOR U4296 ( .A(n4210), .B(n4448), .Z(n4213) );
  XOR U4297 ( .A(n4449), .B(n4450), .Z(n4210) );
  ANDN U4298 ( .A(n4451), .B(n4452), .Z(n4450) );
  XNOR U4299 ( .A(n4449), .B(n4453), .Z(n4451) );
  XOR U4300 ( .A(n4221), .B(n4454), .Z(n4214) );
  IV U4301 ( .A(n4220), .Z(n4454) );
  XNOR U4302 ( .A(n4217), .B(n4455), .Z(n4220) );
  XOR U4303 ( .A(n4456), .B(n4457), .Z(n4217) );
  ANDN U4304 ( .A(n4458), .B(n4459), .Z(n4457) );
  XNOR U4305 ( .A(n4456), .B(n4460), .Z(n4458) );
  XOR U4306 ( .A(n4228), .B(n4461), .Z(n4221) );
  IV U4307 ( .A(n4227), .Z(n4461) );
  XNOR U4308 ( .A(n4224), .B(n4462), .Z(n4227) );
  XOR U4309 ( .A(n4463), .B(n4464), .Z(n4224) );
  ANDN U4310 ( .A(n4465), .B(n4466), .Z(n4464) );
  XNOR U4311 ( .A(n4463), .B(n4467), .Z(n4465) );
  XOR U4312 ( .A(n4235), .B(n4468), .Z(n4228) );
  IV U4313 ( .A(n4234), .Z(n4468) );
  XNOR U4314 ( .A(n4231), .B(n4469), .Z(n4234) );
  XOR U4315 ( .A(n4470), .B(n4471), .Z(n4231) );
  ANDN U4316 ( .A(n4472), .B(n4473), .Z(n4471) );
  XNOR U4317 ( .A(n4470), .B(n4474), .Z(n4472) );
  XOR U4318 ( .A(n4242), .B(n4475), .Z(n4235) );
  IV U4319 ( .A(n4241), .Z(n4475) );
  XNOR U4320 ( .A(n4238), .B(n4476), .Z(n4241) );
  XOR U4321 ( .A(n4477), .B(n4478), .Z(n4238) );
  ANDN U4322 ( .A(n4479), .B(n4480), .Z(n4478) );
  XNOR U4323 ( .A(n4477), .B(n4481), .Z(n4479) );
  XOR U4324 ( .A(n4249), .B(n4482), .Z(n4242) );
  IV U4325 ( .A(n4248), .Z(n4482) );
  XNOR U4326 ( .A(n4245), .B(n4483), .Z(n4248) );
  XOR U4327 ( .A(n4484), .B(n4485), .Z(n4245) );
  ANDN U4328 ( .A(n4486), .B(n4487), .Z(n4485) );
  XNOR U4329 ( .A(n4484), .B(n4488), .Z(n4486) );
  XOR U4330 ( .A(n4256), .B(n4489), .Z(n4249) );
  IV U4331 ( .A(n4255), .Z(n4489) );
  XNOR U4332 ( .A(n4252), .B(n4490), .Z(n4255) );
  XOR U4333 ( .A(n4491), .B(n4492), .Z(n4252) );
  ANDN U4334 ( .A(n4493), .B(n4494), .Z(n4492) );
  XNOR U4335 ( .A(n4491), .B(n4495), .Z(n4493) );
  XOR U4336 ( .A(n4263), .B(n4496), .Z(n4256) );
  IV U4337 ( .A(n4262), .Z(n4496) );
  XNOR U4338 ( .A(n4259), .B(n4497), .Z(n4262) );
  XOR U4339 ( .A(n4498), .B(n4499), .Z(n4259) );
  ANDN U4340 ( .A(n4500), .B(n4501), .Z(n4499) );
  XNOR U4341 ( .A(n4498), .B(n4502), .Z(n4500) );
  XOR U4342 ( .A(n4270), .B(n4503), .Z(n4263) );
  IV U4343 ( .A(n4269), .Z(n4503) );
  XNOR U4344 ( .A(n4266), .B(n4504), .Z(n4269) );
  XOR U4345 ( .A(n4505), .B(n4506), .Z(n4266) );
  ANDN U4346 ( .A(n4507), .B(n4508), .Z(n4506) );
  XNOR U4347 ( .A(n4505), .B(n4509), .Z(n4507) );
  XOR U4348 ( .A(n4277), .B(n4510), .Z(n4270) );
  IV U4349 ( .A(n4276), .Z(n4510) );
  XNOR U4350 ( .A(n4273), .B(n4511), .Z(n4276) );
  XOR U4351 ( .A(n4512), .B(n4513), .Z(n4273) );
  ANDN U4352 ( .A(n4514), .B(n4515), .Z(n4513) );
  XNOR U4353 ( .A(n4512), .B(n4516), .Z(n4514) );
  XOR U4354 ( .A(n4284), .B(n4517), .Z(n4277) );
  IV U4355 ( .A(n4283), .Z(n4517) );
  XNOR U4356 ( .A(n4280), .B(n4518), .Z(n4283) );
  XOR U4357 ( .A(n4519), .B(n4520), .Z(n4280) );
  ANDN U4358 ( .A(n4521), .B(n4522), .Z(n4520) );
  XNOR U4359 ( .A(n4519), .B(n4523), .Z(n4521) );
  XOR U4360 ( .A(n4290), .B(n4524), .Z(n4284) );
  IV U4361 ( .A(n4289), .Z(n4524) );
  XNOR U4362 ( .A(n4286), .B(n4525), .Z(n4289) );
  XOR U4363 ( .A(n4526), .B(n4527), .Z(n4286) );
  ANDN U4364 ( .A(n4528), .B(n4529), .Z(n4527) );
  XNOR U4365 ( .A(n4526), .B(n4530), .Z(n4528) );
  XOR U4366 ( .A(n4296), .B(n4531), .Z(n4290) );
  IV U4367 ( .A(n4295), .Z(n4531) );
  XNOR U4368 ( .A(n4292), .B(n4518), .Z(n4295) );
  AND U4369 ( .A(n5030), .B(n4046), .Z(n4518) );
  XOR U4370 ( .A(n4532), .B(n4533), .Z(n4292) );
  ANDN U4371 ( .A(n4534), .B(n4535), .Z(n4533) );
  XNOR U4372 ( .A(n4532), .B(n4536), .Z(n4534) );
  XOR U4373 ( .A(n4302), .B(n4537), .Z(n4296) );
  IV U4374 ( .A(n4301), .Z(n4537) );
  XNOR U4375 ( .A(n4298), .B(n4511), .Z(n4301) );
  AND U4376 ( .A(n5561), .B(n3593), .Z(n4511) );
  XOR U4377 ( .A(n4538), .B(n4539), .Z(n4298) );
  ANDN U4378 ( .A(n4540), .B(n4541), .Z(n4539) );
  XNOR U4379 ( .A(n4538), .B(n4542), .Z(n4540) );
  XOR U4380 ( .A(n4308), .B(n4543), .Z(n4302) );
  IV U4381 ( .A(n4307), .Z(n4543) );
  XNOR U4382 ( .A(n4304), .B(n4504), .Z(n4307) );
  AND U4383 ( .A(n6118), .B(n3166), .Z(n4504) );
  XOR U4384 ( .A(n4544), .B(n4545), .Z(n4304) );
  ANDN U4385 ( .A(n4546), .B(n4547), .Z(n4545) );
  XNOR U4386 ( .A(n4544), .B(n4548), .Z(n4546) );
  XOR U4387 ( .A(n4314), .B(n4549), .Z(n4308) );
  IV U4388 ( .A(n4313), .Z(n4549) );
  XNOR U4389 ( .A(n4310), .B(n4497), .Z(n4313) );
  AND U4390 ( .A(n6688), .B(n2765), .Z(n4497) );
  XOR U4391 ( .A(n4550), .B(n4551), .Z(n4310) );
  ANDN U4392 ( .A(n4552), .B(n4553), .Z(n4551) );
  XNOR U4393 ( .A(n4550), .B(n4554), .Z(n4552) );
  XOR U4394 ( .A(n4320), .B(n4555), .Z(n4314) );
  IV U4395 ( .A(n4319), .Z(n4555) );
  XNOR U4396 ( .A(n4316), .B(n4490), .Z(n4319) );
  AND U4397 ( .A(n7241), .B(n2396), .Z(n4490) );
  XOR U4398 ( .A(n4556), .B(n4557), .Z(n4316) );
  ANDN U4399 ( .A(n4558), .B(n4559), .Z(n4557) );
  XNOR U4400 ( .A(n4556), .B(n4560), .Z(n4558) );
  XOR U4401 ( .A(n4326), .B(n4561), .Z(n4320) );
  IV U4402 ( .A(n4325), .Z(n4561) );
  XNOR U4403 ( .A(n4322), .B(n4483), .Z(n4325) );
  AND U4404 ( .A(n7770), .B(n2053), .Z(n4483) );
  XOR U4405 ( .A(n4562), .B(n4563), .Z(n4322) );
  ANDN U4406 ( .A(n4564), .B(n4565), .Z(n4563) );
  XNOR U4407 ( .A(n4562), .B(n4566), .Z(n4564) );
  XOR U4408 ( .A(n4332), .B(n4567), .Z(n4326) );
  IV U4409 ( .A(n4331), .Z(n4567) );
  XNOR U4410 ( .A(n4328), .B(n4476), .Z(n4331) );
  AND U4411 ( .A(n8272), .B(n1737), .Z(n4476) );
  XOR U4412 ( .A(n4568), .B(n4569), .Z(n4328) );
  ANDN U4413 ( .A(n4570), .B(n4571), .Z(n4569) );
  XNOR U4414 ( .A(n4568), .B(n4572), .Z(n4570) );
  XOR U4415 ( .A(n4338), .B(n4573), .Z(n4332) );
  IV U4416 ( .A(n4337), .Z(n4573) );
  XNOR U4417 ( .A(n4334), .B(n4469), .Z(n4337) );
  AND U4418 ( .A(n8748), .B(n1448), .Z(n4469) );
  XOR U4419 ( .A(n4574), .B(n4575), .Z(n4334) );
  ANDN U4420 ( .A(n4576), .B(n4577), .Z(n4575) );
  XNOR U4421 ( .A(n4574), .B(n4578), .Z(n4576) );
  XOR U4422 ( .A(n4344), .B(n4579), .Z(n4338) );
  IV U4423 ( .A(n4343), .Z(n4579) );
  XNOR U4424 ( .A(n4340), .B(n4462), .Z(n4343) );
  AND U4425 ( .A(n9198), .B(n1185), .Z(n4462) );
  XOR U4426 ( .A(n4580), .B(n4581), .Z(n4340) );
  ANDN U4427 ( .A(n4582), .B(n4583), .Z(n4581) );
  XNOR U4428 ( .A(n4580), .B(n4584), .Z(n4582) );
  XOR U4429 ( .A(n4350), .B(n4585), .Z(n4344) );
  IV U4430 ( .A(n4349), .Z(n4585) );
  XNOR U4431 ( .A(n4346), .B(n4455), .Z(n4349) );
  AND U4432 ( .A(n9621), .B(n948), .Z(n4455) );
  XOR U4433 ( .A(n4586), .B(n4587), .Z(n4346) );
  ANDN U4434 ( .A(n4588), .B(n4589), .Z(n4587) );
  XNOR U4435 ( .A(n4586), .B(n4590), .Z(n4588) );
  XOR U4436 ( .A(n4356), .B(n4591), .Z(n4350) );
  IV U4437 ( .A(n4355), .Z(n4591) );
  XNOR U4438 ( .A(n4352), .B(n4448), .Z(n4355) );
  AND U4439 ( .A(n10017), .B(n736), .Z(n4448) );
  XOR U4440 ( .A(n4592), .B(n4593), .Z(n4352) );
  ANDN U4441 ( .A(n4594), .B(n4595), .Z(n4593) );
  XNOR U4442 ( .A(n4592), .B(n4596), .Z(n4594) );
  XOR U4443 ( .A(n4362), .B(n4597), .Z(n4356) );
  IV U4444 ( .A(n4361), .Z(n4597) );
  XNOR U4445 ( .A(n4358), .B(n4441), .Z(n4361) );
  AND U4446 ( .A(n10387), .B(n552), .Z(n4441) );
  XOR U4447 ( .A(n4598), .B(n4599), .Z(n4358) );
  ANDN U4448 ( .A(n4600), .B(n4601), .Z(n4599) );
  XNOR U4449 ( .A(n4598), .B(n4602), .Z(n4600) );
  XOR U4450 ( .A(n4368), .B(n4603), .Z(n4362) );
  IV U4451 ( .A(n4367), .Z(n4603) );
  XNOR U4452 ( .A(n4364), .B(n4434), .Z(n4367) );
  AND U4453 ( .A(n10731), .B(n395), .Z(n4434) );
  XOR U4454 ( .A(n4604), .B(n4605), .Z(n4364) );
  ANDN U4455 ( .A(n4606), .B(n4607), .Z(n4605) );
  XNOR U4456 ( .A(n4604), .B(n4608), .Z(n4606) );
  XOR U4457 ( .A(n4374), .B(n4609), .Z(n4368) );
  IV U4458 ( .A(n4373), .Z(n4609) );
  XNOR U4459 ( .A(n4370), .B(n4427), .Z(n4373) );
  AND U4460 ( .A(n11049), .B(n264), .Z(n4427) );
  XOR U4461 ( .A(n4610), .B(n4611), .Z(n4370) );
  ANDN U4462 ( .A(n4612), .B(n4613), .Z(n4611) );
  XNOR U4463 ( .A(n4610), .B(n4614), .Z(n4612) );
  XOR U4464 ( .A(n4380), .B(n4615), .Z(n4374) );
  IV U4465 ( .A(n4379), .Z(n4615) );
  XNOR U4466 ( .A(n4376), .B(n4420), .Z(n4379) );
  AND U4467 ( .A(n11341), .B(n159), .Z(n4420) );
  XOR U4468 ( .A(n4616), .B(n4617), .Z(n4376) );
  ANDN U4469 ( .A(n4618), .B(n4619), .Z(n4617) );
  XNOR U4470 ( .A(n4616), .B(n4620), .Z(n4618) );
  XOR U4471 ( .A(n4387), .B(n4621), .Z(n4380) );
  IV U4472 ( .A(n4386), .Z(n4621) );
  XNOR U4473 ( .A(n4383), .B(n4413), .Z(n4386) );
  AND U4474 ( .A(n11607), .B(n80), .Z(n4413) );
  XOR U4475 ( .A(n4622), .B(n4623), .Z(n4383) );
  ANDN U4476 ( .A(n4624), .B(n4625), .Z(n4623) );
  XNOR U4477 ( .A(n4622), .B(n4626), .Z(n4624) );
  XOR U4478 ( .A(n4392), .B(n4627), .Z(n4387) );
  IV U4479 ( .A(n4391), .Z(n4627) );
  XNOR U4480 ( .A(n4388), .B(n4628), .Z(n4391) );
  AND U4481 ( .A(n42), .B(n11869), .Z(n4628) );
  XOR U4482 ( .A(n4629), .B(n4630), .Z(n4388) );
  ANDN U4483 ( .A(n4631), .B(n4632), .Z(n4630) );
  XNOR U4484 ( .A(n4629), .B(n4633), .Z(n4631) );
  XNOR U4485 ( .A(n4634), .B(n4635), .Z(n4392) );
  ANDN U4486 ( .A(n4636), .B(n4637), .Z(n4635) );
  XNOR U4487 ( .A(n4634), .B(n4638), .Z(n4636) );
  XNOR U4488 ( .A(n4401), .B(n4393), .Z(n4411) );
  XOR U4489 ( .A(n4639), .B(n4640), .Z(n4393) );
  AND U4490 ( .A(n4641), .B(n4642), .Z(n4640) );
  XNOR U4491 ( .A(n4643), .B(n4639), .Z(n4642) );
  XOR U4492 ( .A(n4399), .B(n4644), .Z(n4401) );
  ANDN U4493 ( .A(n11869), .B(n43), .Z(n4644) );
  XOR U4494 ( .A(n4645), .B(n4646), .Z(n4399) );
  AND U4495 ( .A(n4647), .B(n4648), .Z(n4646) );
  XNOR U4496 ( .A(n4645), .B(n4649), .Z(n4648) );
  XOR U4497 ( .A(n4397), .B(n4407), .Z(n4410) );
  XOR U4498 ( .A(n4650), .B(n4651), .Z(n4397) );
  IV U4499 ( .A(n4652), .Z(n4651) );
  XOR U4500 ( .A(n4653), .B(n4654), .Z(n4407) );
  AND U4501 ( .A(n4653), .B(n4655), .Z(n4654) );
  XOR U4502 ( .A(n4656), .B(n4641), .Z(n4655) );
  XOR U4503 ( .A(n4657), .B(n4649), .Z(n4641) );
  XOR U4504 ( .A(n4418), .B(n4658), .Z(n4649) );
  IV U4505 ( .A(n4417), .Z(n4658) );
  XNOR U4506 ( .A(n4414), .B(n4659), .Z(n4417) );
  XOR U4507 ( .A(n4660), .B(n4661), .Z(n4414) );
  ANDN U4508 ( .A(n4662), .B(n4663), .Z(n4661) );
  XNOR U4509 ( .A(n4660), .B(n4664), .Z(n4662) );
  XOR U4510 ( .A(n4425), .B(n4665), .Z(n4418) );
  IV U4511 ( .A(n4424), .Z(n4665) );
  XNOR U4512 ( .A(n4421), .B(n4666), .Z(n4424) );
  XOR U4513 ( .A(n4667), .B(n4668), .Z(n4421) );
  ANDN U4514 ( .A(n4669), .B(n4670), .Z(n4668) );
  XNOR U4515 ( .A(n4667), .B(n4671), .Z(n4669) );
  XOR U4516 ( .A(n4432), .B(n4672), .Z(n4425) );
  IV U4517 ( .A(n4431), .Z(n4672) );
  XNOR U4518 ( .A(n4428), .B(n4673), .Z(n4431) );
  XOR U4519 ( .A(n4674), .B(n4675), .Z(n4428) );
  ANDN U4520 ( .A(n4676), .B(n4677), .Z(n4675) );
  XNOR U4521 ( .A(n4674), .B(n4678), .Z(n4676) );
  XOR U4522 ( .A(n4439), .B(n4679), .Z(n4432) );
  IV U4523 ( .A(n4438), .Z(n4679) );
  XNOR U4524 ( .A(n4435), .B(n4680), .Z(n4438) );
  XOR U4525 ( .A(n4681), .B(n4682), .Z(n4435) );
  ANDN U4526 ( .A(n4683), .B(n4684), .Z(n4682) );
  XNOR U4527 ( .A(n4681), .B(n4685), .Z(n4683) );
  XOR U4528 ( .A(n4446), .B(n4686), .Z(n4439) );
  IV U4529 ( .A(n4445), .Z(n4686) );
  XNOR U4530 ( .A(n4442), .B(n4687), .Z(n4445) );
  XOR U4531 ( .A(n4688), .B(n4689), .Z(n4442) );
  ANDN U4532 ( .A(n4690), .B(n4691), .Z(n4689) );
  XNOR U4533 ( .A(n4688), .B(n4692), .Z(n4690) );
  XOR U4534 ( .A(n4453), .B(n4693), .Z(n4446) );
  IV U4535 ( .A(n4452), .Z(n4693) );
  XNOR U4536 ( .A(n4449), .B(n4694), .Z(n4452) );
  XOR U4537 ( .A(n4695), .B(n4696), .Z(n4449) );
  ANDN U4538 ( .A(n4697), .B(n4698), .Z(n4696) );
  XNOR U4539 ( .A(n4695), .B(n4699), .Z(n4697) );
  XOR U4540 ( .A(n4460), .B(n4700), .Z(n4453) );
  IV U4541 ( .A(n4459), .Z(n4700) );
  XNOR U4542 ( .A(n4456), .B(n4701), .Z(n4459) );
  XOR U4543 ( .A(n4702), .B(n4703), .Z(n4456) );
  ANDN U4544 ( .A(n4704), .B(n4705), .Z(n4703) );
  XNOR U4545 ( .A(n4702), .B(n4706), .Z(n4704) );
  XOR U4546 ( .A(n4467), .B(n4707), .Z(n4460) );
  IV U4547 ( .A(n4466), .Z(n4707) );
  XNOR U4548 ( .A(n4463), .B(n4708), .Z(n4466) );
  XOR U4549 ( .A(n4709), .B(n4710), .Z(n4463) );
  ANDN U4550 ( .A(n4711), .B(n4712), .Z(n4710) );
  XNOR U4551 ( .A(n4709), .B(n4713), .Z(n4711) );
  XOR U4552 ( .A(n4474), .B(n4714), .Z(n4467) );
  IV U4553 ( .A(n4473), .Z(n4714) );
  XNOR U4554 ( .A(n4470), .B(n4715), .Z(n4473) );
  XOR U4555 ( .A(n4716), .B(n4717), .Z(n4470) );
  ANDN U4556 ( .A(n4718), .B(n4719), .Z(n4717) );
  XNOR U4557 ( .A(n4716), .B(n4720), .Z(n4718) );
  XOR U4558 ( .A(n4481), .B(n4721), .Z(n4474) );
  IV U4559 ( .A(n4480), .Z(n4721) );
  XNOR U4560 ( .A(n4477), .B(n4722), .Z(n4480) );
  XOR U4561 ( .A(n4723), .B(n4724), .Z(n4477) );
  ANDN U4562 ( .A(n4725), .B(n4726), .Z(n4724) );
  XNOR U4563 ( .A(n4723), .B(n4727), .Z(n4725) );
  XOR U4564 ( .A(n4488), .B(n4728), .Z(n4481) );
  IV U4565 ( .A(n4487), .Z(n4728) );
  XNOR U4566 ( .A(n4484), .B(n4729), .Z(n4487) );
  XOR U4567 ( .A(n4730), .B(n4731), .Z(n4484) );
  ANDN U4568 ( .A(n4732), .B(n4733), .Z(n4731) );
  XNOR U4569 ( .A(n4730), .B(n4734), .Z(n4732) );
  XOR U4570 ( .A(n4495), .B(n4735), .Z(n4488) );
  IV U4571 ( .A(n4494), .Z(n4735) );
  XNOR U4572 ( .A(n4491), .B(n4736), .Z(n4494) );
  XOR U4573 ( .A(n4737), .B(n4738), .Z(n4491) );
  ANDN U4574 ( .A(n4739), .B(n4740), .Z(n4738) );
  XNOR U4575 ( .A(n4737), .B(n4741), .Z(n4739) );
  XOR U4576 ( .A(n4502), .B(n4742), .Z(n4495) );
  IV U4577 ( .A(n4501), .Z(n4742) );
  XNOR U4578 ( .A(n4498), .B(n4743), .Z(n4501) );
  XOR U4579 ( .A(n4744), .B(n4745), .Z(n4498) );
  ANDN U4580 ( .A(n4746), .B(n4747), .Z(n4745) );
  XNOR U4581 ( .A(n4744), .B(n4748), .Z(n4746) );
  XOR U4582 ( .A(n4509), .B(n4749), .Z(n4502) );
  IV U4583 ( .A(n4508), .Z(n4749) );
  XNOR U4584 ( .A(n4505), .B(n4750), .Z(n4508) );
  XOR U4585 ( .A(n4751), .B(n4752), .Z(n4505) );
  ANDN U4586 ( .A(n4753), .B(n4754), .Z(n4752) );
  XNOR U4587 ( .A(n4751), .B(n4755), .Z(n4753) );
  XOR U4588 ( .A(n4516), .B(n4756), .Z(n4509) );
  IV U4589 ( .A(n4515), .Z(n4756) );
  XNOR U4590 ( .A(n4512), .B(n4757), .Z(n4515) );
  XOR U4591 ( .A(n4758), .B(n4759), .Z(n4512) );
  ANDN U4592 ( .A(n4760), .B(n4761), .Z(n4759) );
  XNOR U4593 ( .A(n4758), .B(n4762), .Z(n4760) );
  XOR U4594 ( .A(n4523), .B(n4763), .Z(n4516) );
  IV U4595 ( .A(n4522), .Z(n4763) );
  XNOR U4596 ( .A(n4519), .B(n4764), .Z(n4522) );
  XOR U4597 ( .A(n4765), .B(n4766), .Z(n4519) );
  ANDN U4598 ( .A(n4767), .B(n4768), .Z(n4766) );
  XNOR U4599 ( .A(n4765), .B(n4769), .Z(n4767) );
  XOR U4600 ( .A(n4530), .B(n4770), .Z(n4523) );
  IV U4601 ( .A(n4529), .Z(n4770) );
  XNOR U4602 ( .A(n4526), .B(n4771), .Z(n4529) );
  XOR U4603 ( .A(n4772), .B(n4773), .Z(n4526) );
  ANDN U4604 ( .A(n4774), .B(n4775), .Z(n4773) );
  XNOR U4605 ( .A(n4772), .B(n4776), .Z(n4774) );
  XOR U4606 ( .A(n4536), .B(n4777), .Z(n4530) );
  IV U4607 ( .A(n4535), .Z(n4777) );
  XNOR U4608 ( .A(n4532), .B(n4771), .Z(n4535) );
  AND U4609 ( .A(n5030), .B(n4525), .Z(n4771) );
  XOR U4610 ( .A(n4778), .B(n4779), .Z(n4532) );
  ANDN U4611 ( .A(n4780), .B(n4781), .Z(n4779) );
  XNOR U4612 ( .A(n4778), .B(n4782), .Z(n4780) );
  XOR U4613 ( .A(n4542), .B(n4783), .Z(n4536) );
  IV U4614 ( .A(n4541), .Z(n4783) );
  XNOR U4615 ( .A(n4538), .B(n4764), .Z(n4541) );
  AND U4616 ( .A(n5561), .B(n4046), .Z(n4764) );
  XOR U4617 ( .A(n4784), .B(n4785), .Z(n4538) );
  ANDN U4618 ( .A(n4786), .B(n4787), .Z(n4785) );
  XNOR U4619 ( .A(n4784), .B(n4788), .Z(n4786) );
  XOR U4620 ( .A(n4548), .B(n4789), .Z(n4542) );
  IV U4621 ( .A(n4547), .Z(n4789) );
  XNOR U4622 ( .A(n4544), .B(n4757), .Z(n4547) );
  AND U4623 ( .A(n6118), .B(n3593), .Z(n4757) );
  XOR U4624 ( .A(n4790), .B(n4791), .Z(n4544) );
  ANDN U4625 ( .A(n4792), .B(n4793), .Z(n4791) );
  XNOR U4626 ( .A(n4790), .B(n4794), .Z(n4792) );
  XOR U4627 ( .A(n4554), .B(n4795), .Z(n4548) );
  IV U4628 ( .A(n4553), .Z(n4795) );
  XNOR U4629 ( .A(n4550), .B(n4750), .Z(n4553) );
  AND U4630 ( .A(n6688), .B(n3166), .Z(n4750) );
  XOR U4631 ( .A(n4796), .B(n4797), .Z(n4550) );
  ANDN U4632 ( .A(n4798), .B(n4799), .Z(n4797) );
  XNOR U4633 ( .A(n4796), .B(n4800), .Z(n4798) );
  XOR U4634 ( .A(n4560), .B(n4801), .Z(n4554) );
  IV U4635 ( .A(n4559), .Z(n4801) );
  XNOR U4636 ( .A(n4556), .B(n4743), .Z(n4559) );
  AND U4637 ( .A(n7241), .B(n2765), .Z(n4743) );
  XOR U4638 ( .A(n4802), .B(n4803), .Z(n4556) );
  ANDN U4639 ( .A(n4804), .B(n4805), .Z(n4803) );
  XNOR U4640 ( .A(n4802), .B(n4806), .Z(n4804) );
  XOR U4641 ( .A(n4566), .B(n4807), .Z(n4560) );
  IV U4642 ( .A(n4565), .Z(n4807) );
  XNOR U4643 ( .A(n4562), .B(n4736), .Z(n4565) );
  AND U4644 ( .A(n7770), .B(n2396), .Z(n4736) );
  XOR U4645 ( .A(n4808), .B(n4809), .Z(n4562) );
  ANDN U4646 ( .A(n4810), .B(n4811), .Z(n4809) );
  XNOR U4647 ( .A(n4808), .B(n4812), .Z(n4810) );
  XOR U4648 ( .A(n4572), .B(n4813), .Z(n4566) );
  IV U4649 ( .A(n4571), .Z(n4813) );
  XNOR U4650 ( .A(n4568), .B(n4729), .Z(n4571) );
  AND U4651 ( .A(n8272), .B(n2053), .Z(n4729) );
  XOR U4652 ( .A(n4814), .B(n4815), .Z(n4568) );
  ANDN U4653 ( .A(n4816), .B(n4817), .Z(n4815) );
  XNOR U4654 ( .A(n4814), .B(n4818), .Z(n4816) );
  XOR U4655 ( .A(n4578), .B(n4819), .Z(n4572) );
  IV U4656 ( .A(n4577), .Z(n4819) );
  XNOR U4657 ( .A(n4574), .B(n4722), .Z(n4577) );
  AND U4658 ( .A(n8748), .B(n1737), .Z(n4722) );
  XOR U4659 ( .A(n4820), .B(n4821), .Z(n4574) );
  ANDN U4660 ( .A(n4822), .B(n4823), .Z(n4821) );
  XNOR U4661 ( .A(n4820), .B(n4824), .Z(n4822) );
  XOR U4662 ( .A(n4584), .B(n4825), .Z(n4578) );
  IV U4663 ( .A(n4583), .Z(n4825) );
  XNOR U4664 ( .A(n4580), .B(n4715), .Z(n4583) );
  AND U4665 ( .A(n9198), .B(n1448), .Z(n4715) );
  XOR U4666 ( .A(n4826), .B(n4827), .Z(n4580) );
  ANDN U4667 ( .A(n4828), .B(n4829), .Z(n4827) );
  XNOR U4668 ( .A(n4826), .B(n4830), .Z(n4828) );
  XOR U4669 ( .A(n4590), .B(n4831), .Z(n4584) );
  IV U4670 ( .A(n4589), .Z(n4831) );
  XNOR U4671 ( .A(n4586), .B(n4708), .Z(n4589) );
  AND U4672 ( .A(n9621), .B(n1185), .Z(n4708) );
  XOR U4673 ( .A(n4832), .B(n4833), .Z(n4586) );
  ANDN U4674 ( .A(n4834), .B(n4835), .Z(n4833) );
  XNOR U4675 ( .A(n4832), .B(n4836), .Z(n4834) );
  XOR U4676 ( .A(n4596), .B(n4837), .Z(n4590) );
  IV U4677 ( .A(n4595), .Z(n4837) );
  XNOR U4678 ( .A(n4592), .B(n4701), .Z(n4595) );
  AND U4679 ( .A(n10017), .B(n948), .Z(n4701) );
  XOR U4680 ( .A(n4838), .B(n4839), .Z(n4592) );
  ANDN U4681 ( .A(n4840), .B(n4841), .Z(n4839) );
  XNOR U4682 ( .A(n4838), .B(n4842), .Z(n4840) );
  XOR U4683 ( .A(n4602), .B(n4843), .Z(n4596) );
  IV U4684 ( .A(n4601), .Z(n4843) );
  XNOR U4685 ( .A(n4598), .B(n4694), .Z(n4601) );
  AND U4686 ( .A(n10387), .B(n736), .Z(n4694) );
  XOR U4687 ( .A(n4844), .B(n4845), .Z(n4598) );
  ANDN U4688 ( .A(n4846), .B(n4847), .Z(n4845) );
  XNOR U4689 ( .A(n4844), .B(n4848), .Z(n4846) );
  XOR U4690 ( .A(n4608), .B(n4849), .Z(n4602) );
  IV U4691 ( .A(n4607), .Z(n4849) );
  XNOR U4692 ( .A(n4604), .B(n4687), .Z(n4607) );
  AND U4693 ( .A(n10731), .B(n552), .Z(n4687) );
  XOR U4694 ( .A(n4850), .B(n4851), .Z(n4604) );
  ANDN U4695 ( .A(n4852), .B(n4853), .Z(n4851) );
  XNOR U4696 ( .A(n4850), .B(n4854), .Z(n4852) );
  XOR U4697 ( .A(n4614), .B(n4855), .Z(n4608) );
  IV U4698 ( .A(n4613), .Z(n4855) );
  XNOR U4699 ( .A(n4610), .B(n4680), .Z(n4613) );
  AND U4700 ( .A(n11049), .B(n395), .Z(n4680) );
  XOR U4701 ( .A(n4856), .B(n4857), .Z(n4610) );
  ANDN U4702 ( .A(n4858), .B(n4859), .Z(n4857) );
  XNOR U4703 ( .A(n4856), .B(n4860), .Z(n4858) );
  XOR U4704 ( .A(n4620), .B(n4861), .Z(n4614) );
  IV U4705 ( .A(n4619), .Z(n4861) );
  XNOR U4706 ( .A(n4616), .B(n4673), .Z(n4619) );
  AND U4707 ( .A(n11341), .B(n264), .Z(n4673) );
  XOR U4708 ( .A(n4862), .B(n4863), .Z(n4616) );
  ANDN U4709 ( .A(n4864), .B(n4865), .Z(n4863) );
  XNOR U4710 ( .A(n4862), .B(n4866), .Z(n4864) );
  XOR U4711 ( .A(n4626), .B(n4867), .Z(n4620) );
  IV U4712 ( .A(n4625), .Z(n4867) );
  XNOR U4713 ( .A(n4622), .B(n4666), .Z(n4625) );
  AND U4714 ( .A(n11607), .B(n159), .Z(n4666) );
  XOR U4715 ( .A(n4868), .B(n4869), .Z(n4622) );
  ANDN U4716 ( .A(n4870), .B(n4871), .Z(n4869) );
  XNOR U4717 ( .A(n4868), .B(n4872), .Z(n4870) );
  XOR U4718 ( .A(n4633), .B(n4873), .Z(n4626) );
  IV U4719 ( .A(n4632), .Z(n4873) );
  XNOR U4720 ( .A(n4629), .B(n4659), .Z(n4632) );
  AND U4721 ( .A(n11869), .B(n80), .Z(n4659) );
  XOR U4722 ( .A(n4874), .B(n4875), .Z(n4629) );
  ANDN U4723 ( .A(n4876), .B(n4877), .Z(n4875) );
  XNOR U4724 ( .A(n4874), .B(n4878), .Z(n4876) );
  XOR U4725 ( .A(n4638), .B(n4879), .Z(n4633) );
  IV U4726 ( .A(n4637), .Z(n4879) );
  XNOR U4727 ( .A(n4634), .B(n4880), .Z(n4637) );
  AND U4728 ( .A(n42), .B(n12128), .Z(n4880) );
  XOR U4729 ( .A(n4881), .B(n4882), .Z(n4634) );
  ANDN U4730 ( .A(n4883), .B(n4884), .Z(n4882) );
  XNOR U4731 ( .A(n4881), .B(n4885), .Z(n4883) );
  XNOR U4732 ( .A(n4886), .B(n4887), .Z(n4638) );
  ANDN U4733 ( .A(n4888), .B(n4889), .Z(n4887) );
  XNOR U4734 ( .A(n4886), .B(n4890), .Z(n4888) );
  XNOR U4735 ( .A(n4647), .B(n4639), .Z(n4657) );
  XOR U4736 ( .A(n4891), .B(n4892), .Z(n4639) );
  AND U4737 ( .A(n4893), .B(n4894), .Z(n4892) );
  XNOR U4738 ( .A(n4895), .B(n4891), .Z(n4894) );
  XOR U4739 ( .A(n4645), .B(n4896), .Z(n4647) );
  ANDN U4740 ( .A(n12128), .B(n43), .Z(n4896) );
  XOR U4741 ( .A(n4897), .B(n4898), .Z(n4645) );
  AND U4742 ( .A(n4899), .B(n4900), .Z(n4898) );
  XNOR U4743 ( .A(n4897), .B(n4901), .Z(n4900) );
  XOR U4744 ( .A(n4643), .B(n4653), .Z(n4656) );
  XOR U4745 ( .A(n4902), .B(n4903), .Z(n4643) );
  IV U4746 ( .A(n4904), .Z(n4903) );
  XOR U4747 ( .A(n4905), .B(n4906), .Z(n4653) );
  AND U4748 ( .A(n4905), .B(n4907), .Z(n4906) );
  XOR U4749 ( .A(n4908), .B(n4893), .Z(n4907) );
  XOR U4750 ( .A(n4909), .B(n4901), .Z(n4893) );
  XOR U4751 ( .A(n4664), .B(n4910), .Z(n4901) );
  IV U4752 ( .A(n4663), .Z(n4910) );
  XNOR U4753 ( .A(n4660), .B(n4911), .Z(n4663) );
  XOR U4754 ( .A(n4912), .B(n4913), .Z(n4660) );
  ANDN U4755 ( .A(n4914), .B(n4915), .Z(n4913) );
  XNOR U4756 ( .A(n4912), .B(n4916), .Z(n4914) );
  XOR U4757 ( .A(n4671), .B(n4917), .Z(n4664) );
  IV U4758 ( .A(n4670), .Z(n4917) );
  XNOR U4759 ( .A(n4667), .B(n4918), .Z(n4670) );
  XOR U4760 ( .A(n4919), .B(n4920), .Z(n4667) );
  ANDN U4761 ( .A(n4921), .B(n4922), .Z(n4920) );
  XNOR U4762 ( .A(n4919), .B(n4923), .Z(n4921) );
  XOR U4763 ( .A(n4678), .B(n4924), .Z(n4671) );
  IV U4764 ( .A(n4677), .Z(n4924) );
  XNOR U4765 ( .A(n4674), .B(n4925), .Z(n4677) );
  XOR U4766 ( .A(n4926), .B(n4927), .Z(n4674) );
  ANDN U4767 ( .A(n4928), .B(n4929), .Z(n4927) );
  XNOR U4768 ( .A(n4926), .B(n4930), .Z(n4928) );
  XOR U4769 ( .A(n4685), .B(n4931), .Z(n4678) );
  IV U4770 ( .A(n4684), .Z(n4931) );
  XNOR U4771 ( .A(n4681), .B(n4932), .Z(n4684) );
  XOR U4772 ( .A(n4933), .B(n4934), .Z(n4681) );
  ANDN U4773 ( .A(n4935), .B(n4936), .Z(n4934) );
  XNOR U4774 ( .A(n4933), .B(n4937), .Z(n4935) );
  XOR U4775 ( .A(n4692), .B(n4938), .Z(n4685) );
  IV U4776 ( .A(n4691), .Z(n4938) );
  XNOR U4777 ( .A(n4688), .B(n4939), .Z(n4691) );
  XOR U4778 ( .A(n4940), .B(n4941), .Z(n4688) );
  ANDN U4779 ( .A(n4942), .B(n4943), .Z(n4941) );
  XNOR U4780 ( .A(n4940), .B(n4944), .Z(n4942) );
  XOR U4781 ( .A(n4699), .B(n4945), .Z(n4692) );
  IV U4782 ( .A(n4698), .Z(n4945) );
  XNOR U4783 ( .A(n4695), .B(n4946), .Z(n4698) );
  XOR U4784 ( .A(n4947), .B(n4948), .Z(n4695) );
  ANDN U4785 ( .A(n4949), .B(n4950), .Z(n4948) );
  XNOR U4786 ( .A(n4947), .B(n4951), .Z(n4949) );
  XOR U4787 ( .A(n4706), .B(n4952), .Z(n4699) );
  IV U4788 ( .A(n4705), .Z(n4952) );
  XNOR U4789 ( .A(n4702), .B(n4953), .Z(n4705) );
  XOR U4790 ( .A(n4954), .B(n4955), .Z(n4702) );
  ANDN U4791 ( .A(n4956), .B(n4957), .Z(n4955) );
  XNOR U4792 ( .A(n4954), .B(n4958), .Z(n4956) );
  XOR U4793 ( .A(n4713), .B(n4959), .Z(n4706) );
  IV U4794 ( .A(n4712), .Z(n4959) );
  XNOR U4795 ( .A(n4709), .B(n4960), .Z(n4712) );
  XOR U4796 ( .A(n4961), .B(n4962), .Z(n4709) );
  ANDN U4797 ( .A(n4963), .B(n4964), .Z(n4962) );
  XNOR U4798 ( .A(n4961), .B(n4965), .Z(n4963) );
  XOR U4799 ( .A(n4720), .B(n4966), .Z(n4713) );
  IV U4800 ( .A(n4719), .Z(n4966) );
  XNOR U4801 ( .A(n4716), .B(n4967), .Z(n4719) );
  XOR U4802 ( .A(n4968), .B(n4969), .Z(n4716) );
  ANDN U4803 ( .A(n4970), .B(n4971), .Z(n4969) );
  XNOR U4804 ( .A(n4968), .B(n4972), .Z(n4970) );
  XOR U4805 ( .A(n4727), .B(n4973), .Z(n4720) );
  IV U4806 ( .A(n4726), .Z(n4973) );
  XNOR U4807 ( .A(n4723), .B(n4974), .Z(n4726) );
  XOR U4808 ( .A(n4975), .B(n4976), .Z(n4723) );
  ANDN U4809 ( .A(n4977), .B(n4978), .Z(n4976) );
  XNOR U4810 ( .A(n4975), .B(n4979), .Z(n4977) );
  XOR U4811 ( .A(n4734), .B(n4980), .Z(n4727) );
  IV U4812 ( .A(n4733), .Z(n4980) );
  XNOR U4813 ( .A(n4730), .B(n4981), .Z(n4733) );
  XOR U4814 ( .A(n4982), .B(n4983), .Z(n4730) );
  ANDN U4815 ( .A(n4984), .B(n4985), .Z(n4983) );
  XNOR U4816 ( .A(n4982), .B(n4986), .Z(n4984) );
  XOR U4817 ( .A(n4741), .B(n4987), .Z(n4734) );
  IV U4818 ( .A(n4740), .Z(n4987) );
  XNOR U4819 ( .A(n4737), .B(n4988), .Z(n4740) );
  XOR U4820 ( .A(n4989), .B(n4990), .Z(n4737) );
  ANDN U4821 ( .A(n4991), .B(n4992), .Z(n4990) );
  XNOR U4822 ( .A(n4989), .B(n4993), .Z(n4991) );
  XOR U4823 ( .A(n4748), .B(n4994), .Z(n4741) );
  IV U4824 ( .A(n4747), .Z(n4994) );
  XNOR U4825 ( .A(n4744), .B(n4995), .Z(n4747) );
  XOR U4826 ( .A(n4996), .B(n4997), .Z(n4744) );
  ANDN U4827 ( .A(n4998), .B(n4999), .Z(n4997) );
  XNOR U4828 ( .A(n4996), .B(n5000), .Z(n4998) );
  XOR U4829 ( .A(n4755), .B(n5001), .Z(n4748) );
  IV U4830 ( .A(n4754), .Z(n5001) );
  XNOR U4831 ( .A(n4751), .B(n5002), .Z(n4754) );
  XOR U4832 ( .A(n5003), .B(n5004), .Z(n4751) );
  ANDN U4833 ( .A(n5005), .B(n5006), .Z(n5004) );
  XNOR U4834 ( .A(n5003), .B(n5007), .Z(n5005) );
  XOR U4835 ( .A(n4762), .B(n5008), .Z(n4755) );
  IV U4836 ( .A(n4761), .Z(n5008) );
  XNOR U4837 ( .A(n4758), .B(n5009), .Z(n4761) );
  XOR U4838 ( .A(n5010), .B(n5011), .Z(n4758) );
  ANDN U4839 ( .A(n5012), .B(n5013), .Z(n5011) );
  XNOR U4840 ( .A(n5010), .B(n5014), .Z(n5012) );
  XOR U4841 ( .A(n4769), .B(n5015), .Z(n4762) );
  IV U4842 ( .A(n4768), .Z(n5015) );
  XNOR U4843 ( .A(n4765), .B(n5016), .Z(n4768) );
  XOR U4844 ( .A(n5017), .B(n5018), .Z(n4765) );
  ANDN U4845 ( .A(n5019), .B(n5020), .Z(n5018) );
  XNOR U4846 ( .A(n5017), .B(n5021), .Z(n5019) );
  XOR U4847 ( .A(n4776), .B(n5022), .Z(n4769) );
  IV U4848 ( .A(n4775), .Z(n5022) );
  XNOR U4849 ( .A(n4772), .B(n5023), .Z(n4775) );
  XOR U4850 ( .A(n5024), .B(n5025), .Z(n4772) );
  ANDN U4851 ( .A(n5026), .B(n5027), .Z(n5025) );
  XNOR U4852 ( .A(n5024), .B(n5028), .Z(n5026) );
  XOR U4853 ( .A(n4782), .B(n5029), .Z(n4776) );
  IV U4854 ( .A(n4781), .Z(n5029) );
  XNOR U4855 ( .A(n4778), .B(n5030), .Z(n4781) );
  XOR U4856 ( .A(n5031), .B(n5032), .Z(n4778) );
  ANDN U4857 ( .A(n5033), .B(n5034), .Z(n5032) );
  XNOR U4858 ( .A(n5031), .B(n5035), .Z(n5033) );
  XOR U4859 ( .A(n4788), .B(n5036), .Z(n4782) );
  IV U4860 ( .A(n4787), .Z(n5036) );
  XNOR U4861 ( .A(n4784), .B(n5023), .Z(n4787) );
  AND U4862 ( .A(n5561), .B(n4525), .Z(n5023) );
  XOR U4863 ( .A(n5037), .B(n5038), .Z(n4784) );
  ANDN U4864 ( .A(n5039), .B(n5040), .Z(n5038) );
  XNOR U4865 ( .A(n5037), .B(n5041), .Z(n5039) );
  XOR U4866 ( .A(n4794), .B(n5042), .Z(n4788) );
  IV U4867 ( .A(n4793), .Z(n5042) );
  XNOR U4868 ( .A(n4790), .B(n5016), .Z(n4793) );
  AND U4869 ( .A(n6118), .B(n4046), .Z(n5016) );
  XOR U4870 ( .A(n5043), .B(n5044), .Z(n4790) );
  ANDN U4871 ( .A(n5045), .B(n5046), .Z(n5044) );
  XNOR U4872 ( .A(n5043), .B(n5047), .Z(n5045) );
  XOR U4873 ( .A(n4800), .B(n5048), .Z(n4794) );
  IV U4874 ( .A(n4799), .Z(n5048) );
  XNOR U4875 ( .A(n4796), .B(n5009), .Z(n4799) );
  AND U4876 ( .A(n6688), .B(n3593), .Z(n5009) );
  XOR U4877 ( .A(n5049), .B(n5050), .Z(n4796) );
  ANDN U4878 ( .A(n5051), .B(n5052), .Z(n5050) );
  XNOR U4879 ( .A(n5049), .B(n5053), .Z(n5051) );
  XOR U4880 ( .A(n4806), .B(n5054), .Z(n4800) );
  IV U4881 ( .A(n4805), .Z(n5054) );
  XNOR U4882 ( .A(n4802), .B(n5002), .Z(n4805) );
  AND U4883 ( .A(n7241), .B(n3166), .Z(n5002) );
  XOR U4884 ( .A(n5055), .B(n5056), .Z(n4802) );
  ANDN U4885 ( .A(n5057), .B(n5058), .Z(n5056) );
  XNOR U4886 ( .A(n5055), .B(n5059), .Z(n5057) );
  XOR U4887 ( .A(n4812), .B(n5060), .Z(n4806) );
  IV U4888 ( .A(n4811), .Z(n5060) );
  XNOR U4889 ( .A(n4808), .B(n4995), .Z(n4811) );
  AND U4890 ( .A(n7770), .B(n2765), .Z(n4995) );
  XOR U4891 ( .A(n5061), .B(n5062), .Z(n4808) );
  ANDN U4892 ( .A(n5063), .B(n5064), .Z(n5062) );
  XNOR U4893 ( .A(n5061), .B(n5065), .Z(n5063) );
  XOR U4894 ( .A(n4818), .B(n5066), .Z(n4812) );
  IV U4895 ( .A(n4817), .Z(n5066) );
  XNOR U4896 ( .A(n4814), .B(n4988), .Z(n4817) );
  AND U4897 ( .A(n8272), .B(n2396), .Z(n4988) );
  XOR U4898 ( .A(n5067), .B(n5068), .Z(n4814) );
  ANDN U4899 ( .A(n5069), .B(n5070), .Z(n5068) );
  XNOR U4900 ( .A(n5067), .B(n5071), .Z(n5069) );
  XOR U4901 ( .A(n4824), .B(n5072), .Z(n4818) );
  IV U4902 ( .A(n4823), .Z(n5072) );
  XNOR U4903 ( .A(n4820), .B(n4981), .Z(n4823) );
  AND U4904 ( .A(n8748), .B(n2053), .Z(n4981) );
  XOR U4905 ( .A(n5073), .B(n5074), .Z(n4820) );
  ANDN U4906 ( .A(n5075), .B(n5076), .Z(n5074) );
  XNOR U4907 ( .A(n5073), .B(n5077), .Z(n5075) );
  XOR U4908 ( .A(n4830), .B(n5078), .Z(n4824) );
  IV U4909 ( .A(n4829), .Z(n5078) );
  XNOR U4910 ( .A(n4826), .B(n4974), .Z(n4829) );
  AND U4911 ( .A(n9198), .B(n1737), .Z(n4974) );
  XOR U4912 ( .A(n5079), .B(n5080), .Z(n4826) );
  ANDN U4913 ( .A(n5081), .B(n5082), .Z(n5080) );
  XNOR U4914 ( .A(n5079), .B(n5083), .Z(n5081) );
  XOR U4915 ( .A(n4836), .B(n5084), .Z(n4830) );
  IV U4916 ( .A(n4835), .Z(n5084) );
  XNOR U4917 ( .A(n4832), .B(n4967), .Z(n4835) );
  AND U4918 ( .A(n9621), .B(n1448), .Z(n4967) );
  XOR U4919 ( .A(n5085), .B(n5086), .Z(n4832) );
  ANDN U4920 ( .A(n5087), .B(n5088), .Z(n5086) );
  XNOR U4921 ( .A(n5085), .B(n5089), .Z(n5087) );
  XOR U4922 ( .A(n4842), .B(n5090), .Z(n4836) );
  IV U4923 ( .A(n4841), .Z(n5090) );
  XNOR U4924 ( .A(n4838), .B(n4960), .Z(n4841) );
  AND U4925 ( .A(n10017), .B(n1185), .Z(n4960) );
  XOR U4926 ( .A(n5091), .B(n5092), .Z(n4838) );
  ANDN U4927 ( .A(n5093), .B(n5094), .Z(n5092) );
  XNOR U4928 ( .A(n5091), .B(n5095), .Z(n5093) );
  XOR U4929 ( .A(n4848), .B(n5096), .Z(n4842) );
  IV U4930 ( .A(n4847), .Z(n5096) );
  XNOR U4931 ( .A(n4844), .B(n4953), .Z(n4847) );
  AND U4932 ( .A(n10387), .B(n948), .Z(n4953) );
  XOR U4933 ( .A(n5097), .B(n5098), .Z(n4844) );
  ANDN U4934 ( .A(n5099), .B(n5100), .Z(n5098) );
  XNOR U4935 ( .A(n5097), .B(n5101), .Z(n5099) );
  XOR U4936 ( .A(n4854), .B(n5102), .Z(n4848) );
  IV U4937 ( .A(n4853), .Z(n5102) );
  XNOR U4938 ( .A(n4850), .B(n4946), .Z(n4853) );
  AND U4939 ( .A(n10731), .B(n736), .Z(n4946) );
  XOR U4940 ( .A(n5103), .B(n5104), .Z(n4850) );
  ANDN U4941 ( .A(n5105), .B(n5106), .Z(n5104) );
  XNOR U4942 ( .A(n5103), .B(n5107), .Z(n5105) );
  XOR U4943 ( .A(n4860), .B(n5108), .Z(n4854) );
  IV U4944 ( .A(n4859), .Z(n5108) );
  XNOR U4945 ( .A(n4856), .B(n4939), .Z(n4859) );
  AND U4946 ( .A(n11049), .B(n552), .Z(n4939) );
  XOR U4947 ( .A(n5109), .B(n5110), .Z(n4856) );
  ANDN U4948 ( .A(n5111), .B(n5112), .Z(n5110) );
  XNOR U4949 ( .A(n5109), .B(n5113), .Z(n5111) );
  XOR U4950 ( .A(n4866), .B(n5114), .Z(n4860) );
  IV U4951 ( .A(n4865), .Z(n5114) );
  XNOR U4952 ( .A(n4862), .B(n4932), .Z(n4865) );
  AND U4953 ( .A(n11341), .B(n395), .Z(n4932) );
  XOR U4954 ( .A(n5115), .B(n5116), .Z(n4862) );
  ANDN U4955 ( .A(n5117), .B(n5118), .Z(n5116) );
  XNOR U4956 ( .A(n5115), .B(n5119), .Z(n5117) );
  XOR U4957 ( .A(n4872), .B(n5120), .Z(n4866) );
  IV U4958 ( .A(n4871), .Z(n5120) );
  XNOR U4959 ( .A(n4868), .B(n4925), .Z(n4871) );
  AND U4960 ( .A(n11607), .B(n264), .Z(n4925) );
  XOR U4961 ( .A(n5121), .B(n5122), .Z(n4868) );
  ANDN U4962 ( .A(n5123), .B(n5124), .Z(n5122) );
  XNOR U4963 ( .A(n5121), .B(n5125), .Z(n5123) );
  XOR U4964 ( .A(n4878), .B(n5126), .Z(n4872) );
  IV U4965 ( .A(n4877), .Z(n5126) );
  XNOR U4966 ( .A(n4874), .B(n4918), .Z(n4877) );
  AND U4967 ( .A(n11869), .B(n159), .Z(n4918) );
  XOR U4968 ( .A(n5127), .B(n5128), .Z(n4874) );
  ANDN U4969 ( .A(n5129), .B(n5130), .Z(n5128) );
  XNOR U4970 ( .A(n5127), .B(n5131), .Z(n5129) );
  XOR U4971 ( .A(n4885), .B(n5132), .Z(n4878) );
  IV U4972 ( .A(n4884), .Z(n5132) );
  XNOR U4973 ( .A(n4881), .B(n4911), .Z(n4884) );
  AND U4974 ( .A(n12128), .B(n80), .Z(n4911) );
  XOR U4975 ( .A(n5133), .B(n5134), .Z(n4881) );
  ANDN U4976 ( .A(n5135), .B(n5136), .Z(n5134) );
  XNOR U4977 ( .A(n5133), .B(n5137), .Z(n5135) );
  XOR U4978 ( .A(n4890), .B(n5138), .Z(n4885) );
  IV U4979 ( .A(n4889), .Z(n5138) );
  XNOR U4980 ( .A(n4886), .B(n5139), .Z(n4889) );
  AND U4981 ( .A(n42), .B(n12387), .Z(n5139) );
  XOR U4982 ( .A(n5140), .B(n5141), .Z(n4886) );
  ANDN U4983 ( .A(n5142), .B(n5143), .Z(n5141) );
  XNOR U4984 ( .A(n5140), .B(n5144), .Z(n5142) );
  XNOR U4985 ( .A(n5145), .B(n5146), .Z(n4890) );
  ANDN U4986 ( .A(n5147), .B(n5148), .Z(n5146) );
  XNOR U4987 ( .A(n5145), .B(n5149), .Z(n5147) );
  XNOR U4988 ( .A(n4899), .B(n4891), .Z(n4909) );
  XOR U4989 ( .A(n5150), .B(n5151), .Z(n4891) );
  AND U4990 ( .A(n5152), .B(n5153), .Z(n5151) );
  XNOR U4991 ( .A(n5154), .B(n5150), .Z(n5153) );
  XOR U4992 ( .A(n4897), .B(n5155), .Z(n4899) );
  ANDN U4993 ( .A(n12387), .B(n43), .Z(n5155) );
  XOR U4994 ( .A(n5156), .B(n5157), .Z(n4897) );
  AND U4995 ( .A(n5158), .B(n5159), .Z(n5157) );
  XNOR U4996 ( .A(n5156), .B(n5160), .Z(n5159) );
  XOR U4997 ( .A(n4895), .B(n4905), .Z(n4908) );
  XOR U4998 ( .A(n5161), .B(n5162), .Z(n4895) );
  IV U4999 ( .A(n5163), .Z(n5162) );
  XOR U5000 ( .A(n5164), .B(n5165), .Z(n4905) );
  AND U5001 ( .A(n5164), .B(n5166), .Z(n5165) );
  XOR U5002 ( .A(n5167), .B(n5152), .Z(n5166) );
  XOR U5003 ( .A(n5168), .B(n5160), .Z(n5152) );
  XOR U5004 ( .A(n4916), .B(n5169), .Z(n5160) );
  IV U5005 ( .A(n4915), .Z(n5169) );
  XNOR U5006 ( .A(n4912), .B(n5170), .Z(n4915) );
  XOR U5007 ( .A(n5171), .B(n5172), .Z(n4912) );
  ANDN U5008 ( .A(n5173), .B(n5174), .Z(n5172) );
  XNOR U5009 ( .A(n5171), .B(n5175), .Z(n5173) );
  XOR U5010 ( .A(n4923), .B(n5176), .Z(n4916) );
  IV U5011 ( .A(n4922), .Z(n5176) );
  XNOR U5012 ( .A(n4919), .B(n5177), .Z(n4922) );
  XOR U5013 ( .A(n5178), .B(n5179), .Z(n4919) );
  ANDN U5014 ( .A(n5180), .B(n5181), .Z(n5179) );
  XNOR U5015 ( .A(n5178), .B(n5182), .Z(n5180) );
  XOR U5016 ( .A(n4930), .B(n5183), .Z(n4923) );
  IV U5017 ( .A(n4929), .Z(n5183) );
  XNOR U5018 ( .A(n4926), .B(n5184), .Z(n4929) );
  XOR U5019 ( .A(n5185), .B(n5186), .Z(n4926) );
  ANDN U5020 ( .A(n5187), .B(n5188), .Z(n5186) );
  XNOR U5021 ( .A(n5185), .B(n5189), .Z(n5187) );
  XOR U5022 ( .A(n4937), .B(n5190), .Z(n4930) );
  IV U5023 ( .A(n4936), .Z(n5190) );
  XNOR U5024 ( .A(n4933), .B(n5191), .Z(n4936) );
  XOR U5025 ( .A(n5192), .B(n5193), .Z(n4933) );
  ANDN U5026 ( .A(n5194), .B(n5195), .Z(n5193) );
  XNOR U5027 ( .A(n5192), .B(n5196), .Z(n5194) );
  XOR U5028 ( .A(n4944), .B(n5197), .Z(n4937) );
  IV U5029 ( .A(n4943), .Z(n5197) );
  XNOR U5030 ( .A(n4940), .B(n5198), .Z(n4943) );
  XOR U5031 ( .A(n5199), .B(n5200), .Z(n4940) );
  ANDN U5032 ( .A(n5201), .B(n5202), .Z(n5200) );
  XNOR U5033 ( .A(n5199), .B(n5203), .Z(n5201) );
  XOR U5034 ( .A(n4951), .B(n5204), .Z(n4944) );
  IV U5035 ( .A(n4950), .Z(n5204) );
  XNOR U5036 ( .A(n4947), .B(n5205), .Z(n4950) );
  XOR U5037 ( .A(n5206), .B(n5207), .Z(n4947) );
  ANDN U5038 ( .A(n5208), .B(n5209), .Z(n5207) );
  XNOR U5039 ( .A(n5206), .B(n5210), .Z(n5208) );
  XOR U5040 ( .A(n4958), .B(n5211), .Z(n4951) );
  IV U5041 ( .A(n4957), .Z(n5211) );
  XNOR U5042 ( .A(n4954), .B(n5212), .Z(n4957) );
  XOR U5043 ( .A(n5213), .B(n5214), .Z(n4954) );
  ANDN U5044 ( .A(n5215), .B(n5216), .Z(n5214) );
  XNOR U5045 ( .A(n5213), .B(n5217), .Z(n5215) );
  XOR U5046 ( .A(n4965), .B(n5218), .Z(n4958) );
  IV U5047 ( .A(n4964), .Z(n5218) );
  XNOR U5048 ( .A(n4961), .B(n5219), .Z(n4964) );
  XOR U5049 ( .A(n5220), .B(n5221), .Z(n4961) );
  ANDN U5050 ( .A(n5222), .B(n5223), .Z(n5221) );
  XNOR U5051 ( .A(n5220), .B(n5224), .Z(n5222) );
  XOR U5052 ( .A(n4972), .B(n5225), .Z(n4965) );
  IV U5053 ( .A(n4971), .Z(n5225) );
  XNOR U5054 ( .A(n4968), .B(n5226), .Z(n4971) );
  XOR U5055 ( .A(n5227), .B(n5228), .Z(n4968) );
  ANDN U5056 ( .A(n5229), .B(n5230), .Z(n5228) );
  XNOR U5057 ( .A(n5227), .B(n5231), .Z(n5229) );
  XOR U5058 ( .A(n4979), .B(n5232), .Z(n4972) );
  IV U5059 ( .A(n4978), .Z(n5232) );
  XNOR U5060 ( .A(n4975), .B(n5233), .Z(n4978) );
  XOR U5061 ( .A(n5234), .B(n5235), .Z(n4975) );
  ANDN U5062 ( .A(n5236), .B(n5237), .Z(n5235) );
  XNOR U5063 ( .A(n5234), .B(n5238), .Z(n5236) );
  XOR U5064 ( .A(n4986), .B(n5239), .Z(n4979) );
  IV U5065 ( .A(n4985), .Z(n5239) );
  XNOR U5066 ( .A(n4982), .B(n5240), .Z(n4985) );
  XOR U5067 ( .A(n5241), .B(n5242), .Z(n4982) );
  ANDN U5068 ( .A(n5243), .B(n5244), .Z(n5242) );
  XNOR U5069 ( .A(n5241), .B(n5245), .Z(n5243) );
  XOR U5070 ( .A(n4993), .B(n5246), .Z(n4986) );
  IV U5071 ( .A(n4992), .Z(n5246) );
  XNOR U5072 ( .A(n4989), .B(n5247), .Z(n4992) );
  XOR U5073 ( .A(n5248), .B(n5249), .Z(n4989) );
  ANDN U5074 ( .A(n5250), .B(n5251), .Z(n5249) );
  XNOR U5075 ( .A(n5248), .B(n5252), .Z(n5250) );
  XOR U5076 ( .A(n5000), .B(n5253), .Z(n4993) );
  IV U5077 ( .A(n4999), .Z(n5253) );
  XNOR U5078 ( .A(n4996), .B(n5254), .Z(n4999) );
  XOR U5079 ( .A(n5255), .B(n5256), .Z(n4996) );
  ANDN U5080 ( .A(n5257), .B(n5258), .Z(n5256) );
  XNOR U5081 ( .A(n5255), .B(n5259), .Z(n5257) );
  XOR U5082 ( .A(n5007), .B(n5260), .Z(n5000) );
  IV U5083 ( .A(n5006), .Z(n5260) );
  XNOR U5084 ( .A(n5003), .B(n5261), .Z(n5006) );
  XOR U5085 ( .A(n5262), .B(n5263), .Z(n5003) );
  ANDN U5086 ( .A(n5264), .B(n5265), .Z(n5263) );
  XNOR U5087 ( .A(n5262), .B(n5266), .Z(n5264) );
  XOR U5088 ( .A(n5014), .B(n5267), .Z(n5007) );
  IV U5089 ( .A(n5013), .Z(n5267) );
  XNOR U5090 ( .A(n5010), .B(n5268), .Z(n5013) );
  XOR U5091 ( .A(n5269), .B(n5270), .Z(n5010) );
  ANDN U5092 ( .A(n5271), .B(n5272), .Z(n5270) );
  XNOR U5093 ( .A(n5269), .B(n5273), .Z(n5271) );
  XOR U5094 ( .A(n5021), .B(n5274), .Z(n5014) );
  IV U5095 ( .A(n5020), .Z(n5274) );
  XNOR U5096 ( .A(n5017), .B(n5275), .Z(n5020) );
  XOR U5097 ( .A(n5276), .B(n5277), .Z(n5017) );
  ANDN U5098 ( .A(n5278), .B(n5279), .Z(n5277) );
  XNOR U5099 ( .A(n5276), .B(n5280), .Z(n5278) );
  XOR U5100 ( .A(n5028), .B(n5281), .Z(n5021) );
  IV U5101 ( .A(n5027), .Z(n5281) );
  XNOR U5102 ( .A(n5024), .B(n5282), .Z(n5027) );
  XOR U5103 ( .A(n5283), .B(n5284), .Z(n5024) );
  ANDN U5104 ( .A(n5285), .B(n5286), .Z(n5284) );
  XNOR U5105 ( .A(n5283), .B(n5287), .Z(n5285) );
  XOR U5106 ( .A(n5035), .B(n5288), .Z(n5028) );
  IV U5107 ( .A(n5034), .Z(n5288) );
  XNOR U5108 ( .A(n5031), .B(n5289), .Z(n5034) );
  XOR U5109 ( .A(n5290), .B(n5291), .Z(n5031) );
  ANDN U5110 ( .A(n5292), .B(n5293), .Z(n5291) );
  XNOR U5111 ( .A(n5290), .B(n5294), .Z(n5292) );
  XOR U5112 ( .A(n5041), .B(n5295), .Z(n5035) );
  IV U5113 ( .A(n5040), .Z(n5295) );
  XNOR U5114 ( .A(n5037), .B(n5289), .Z(n5040) );
  AND U5115 ( .A(n5561), .B(n5030), .Z(n5289) );
  XOR U5116 ( .A(n5296), .B(n5297), .Z(n5037) );
  ANDN U5117 ( .A(n5298), .B(n5299), .Z(n5297) );
  XNOR U5118 ( .A(n5296), .B(n5300), .Z(n5298) );
  XOR U5119 ( .A(n5047), .B(n5301), .Z(n5041) );
  IV U5120 ( .A(n5046), .Z(n5301) );
  XNOR U5121 ( .A(n5043), .B(n5282), .Z(n5046) );
  AND U5122 ( .A(n6118), .B(n4525), .Z(n5282) );
  XOR U5123 ( .A(n5302), .B(n5303), .Z(n5043) );
  ANDN U5124 ( .A(n5304), .B(n5305), .Z(n5303) );
  XNOR U5125 ( .A(n5302), .B(n5306), .Z(n5304) );
  XOR U5126 ( .A(n5053), .B(n5307), .Z(n5047) );
  IV U5127 ( .A(n5052), .Z(n5307) );
  XNOR U5128 ( .A(n5049), .B(n5275), .Z(n5052) );
  AND U5129 ( .A(n6688), .B(n4046), .Z(n5275) );
  XOR U5130 ( .A(n5308), .B(n5309), .Z(n5049) );
  ANDN U5131 ( .A(n5310), .B(n5311), .Z(n5309) );
  XNOR U5132 ( .A(n5308), .B(n5312), .Z(n5310) );
  XOR U5133 ( .A(n5059), .B(n5313), .Z(n5053) );
  IV U5134 ( .A(n5058), .Z(n5313) );
  XNOR U5135 ( .A(n5055), .B(n5268), .Z(n5058) );
  AND U5136 ( .A(n7241), .B(n3593), .Z(n5268) );
  XOR U5137 ( .A(n5314), .B(n5315), .Z(n5055) );
  ANDN U5138 ( .A(n5316), .B(n5317), .Z(n5315) );
  XNOR U5139 ( .A(n5314), .B(n5318), .Z(n5316) );
  XOR U5140 ( .A(n5065), .B(n5319), .Z(n5059) );
  IV U5141 ( .A(n5064), .Z(n5319) );
  XNOR U5142 ( .A(n5061), .B(n5261), .Z(n5064) );
  AND U5143 ( .A(n7770), .B(n3166), .Z(n5261) );
  XOR U5144 ( .A(n5320), .B(n5321), .Z(n5061) );
  ANDN U5145 ( .A(n5322), .B(n5323), .Z(n5321) );
  XNOR U5146 ( .A(n5320), .B(n5324), .Z(n5322) );
  XOR U5147 ( .A(n5071), .B(n5325), .Z(n5065) );
  IV U5148 ( .A(n5070), .Z(n5325) );
  XNOR U5149 ( .A(n5067), .B(n5254), .Z(n5070) );
  AND U5150 ( .A(n8272), .B(n2765), .Z(n5254) );
  XOR U5151 ( .A(n5326), .B(n5327), .Z(n5067) );
  ANDN U5152 ( .A(n5328), .B(n5329), .Z(n5327) );
  XNOR U5153 ( .A(n5326), .B(n5330), .Z(n5328) );
  XOR U5154 ( .A(n5077), .B(n5331), .Z(n5071) );
  IV U5155 ( .A(n5076), .Z(n5331) );
  XNOR U5156 ( .A(n5073), .B(n5247), .Z(n5076) );
  AND U5157 ( .A(n8748), .B(n2396), .Z(n5247) );
  XOR U5158 ( .A(n5332), .B(n5333), .Z(n5073) );
  ANDN U5159 ( .A(n5334), .B(n5335), .Z(n5333) );
  XNOR U5160 ( .A(n5332), .B(n5336), .Z(n5334) );
  XOR U5161 ( .A(n5083), .B(n5337), .Z(n5077) );
  IV U5162 ( .A(n5082), .Z(n5337) );
  XNOR U5163 ( .A(n5079), .B(n5240), .Z(n5082) );
  AND U5164 ( .A(n9198), .B(n2053), .Z(n5240) );
  XOR U5165 ( .A(n5338), .B(n5339), .Z(n5079) );
  ANDN U5166 ( .A(n5340), .B(n5341), .Z(n5339) );
  XNOR U5167 ( .A(n5338), .B(n5342), .Z(n5340) );
  XOR U5168 ( .A(n5089), .B(n5343), .Z(n5083) );
  IV U5169 ( .A(n5088), .Z(n5343) );
  XNOR U5170 ( .A(n5085), .B(n5233), .Z(n5088) );
  AND U5171 ( .A(n9621), .B(n1737), .Z(n5233) );
  XOR U5172 ( .A(n5344), .B(n5345), .Z(n5085) );
  ANDN U5173 ( .A(n5346), .B(n5347), .Z(n5345) );
  XNOR U5174 ( .A(n5344), .B(n5348), .Z(n5346) );
  XOR U5175 ( .A(n5095), .B(n5349), .Z(n5089) );
  IV U5176 ( .A(n5094), .Z(n5349) );
  XNOR U5177 ( .A(n5091), .B(n5226), .Z(n5094) );
  AND U5178 ( .A(n10017), .B(n1448), .Z(n5226) );
  XOR U5179 ( .A(n5350), .B(n5351), .Z(n5091) );
  ANDN U5180 ( .A(n5352), .B(n5353), .Z(n5351) );
  XNOR U5181 ( .A(n5350), .B(n5354), .Z(n5352) );
  XOR U5182 ( .A(n5101), .B(n5355), .Z(n5095) );
  IV U5183 ( .A(n5100), .Z(n5355) );
  XNOR U5184 ( .A(n5097), .B(n5219), .Z(n5100) );
  AND U5185 ( .A(n10387), .B(n1185), .Z(n5219) );
  XOR U5186 ( .A(n5356), .B(n5357), .Z(n5097) );
  ANDN U5187 ( .A(n5358), .B(n5359), .Z(n5357) );
  XNOR U5188 ( .A(n5356), .B(n5360), .Z(n5358) );
  XOR U5189 ( .A(n5107), .B(n5361), .Z(n5101) );
  IV U5190 ( .A(n5106), .Z(n5361) );
  XNOR U5191 ( .A(n5103), .B(n5212), .Z(n5106) );
  AND U5192 ( .A(n10731), .B(n948), .Z(n5212) );
  XOR U5193 ( .A(n5362), .B(n5363), .Z(n5103) );
  ANDN U5194 ( .A(n5364), .B(n5365), .Z(n5363) );
  XNOR U5195 ( .A(n5362), .B(n5366), .Z(n5364) );
  XOR U5196 ( .A(n5113), .B(n5367), .Z(n5107) );
  IV U5197 ( .A(n5112), .Z(n5367) );
  XNOR U5198 ( .A(n5109), .B(n5205), .Z(n5112) );
  AND U5199 ( .A(n11049), .B(n736), .Z(n5205) );
  XOR U5200 ( .A(n5368), .B(n5369), .Z(n5109) );
  ANDN U5201 ( .A(n5370), .B(n5371), .Z(n5369) );
  XNOR U5202 ( .A(n5368), .B(n5372), .Z(n5370) );
  XOR U5203 ( .A(n5119), .B(n5373), .Z(n5113) );
  IV U5204 ( .A(n5118), .Z(n5373) );
  XNOR U5205 ( .A(n5115), .B(n5198), .Z(n5118) );
  AND U5206 ( .A(n11341), .B(n552), .Z(n5198) );
  XOR U5207 ( .A(n5374), .B(n5375), .Z(n5115) );
  ANDN U5208 ( .A(n5376), .B(n5377), .Z(n5375) );
  XNOR U5209 ( .A(n5374), .B(n5378), .Z(n5376) );
  XOR U5210 ( .A(n5125), .B(n5379), .Z(n5119) );
  IV U5211 ( .A(n5124), .Z(n5379) );
  XNOR U5212 ( .A(n5121), .B(n5191), .Z(n5124) );
  AND U5213 ( .A(n11607), .B(n395), .Z(n5191) );
  XOR U5214 ( .A(n5380), .B(n5381), .Z(n5121) );
  ANDN U5215 ( .A(n5382), .B(n5383), .Z(n5381) );
  XNOR U5216 ( .A(n5380), .B(n5384), .Z(n5382) );
  XOR U5217 ( .A(n5131), .B(n5385), .Z(n5125) );
  IV U5218 ( .A(n5130), .Z(n5385) );
  XNOR U5219 ( .A(n5127), .B(n5184), .Z(n5130) );
  AND U5220 ( .A(n11869), .B(n264), .Z(n5184) );
  XOR U5221 ( .A(n5386), .B(n5387), .Z(n5127) );
  ANDN U5222 ( .A(n5388), .B(n5389), .Z(n5387) );
  XNOR U5223 ( .A(n5386), .B(n5390), .Z(n5388) );
  XOR U5224 ( .A(n5137), .B(n5391), .Z(n5131) );
  IV U5225 ( .A(n5136), .Z(n5391) );
  XNOR U5226 ( .A(n5133), .B(n5177), .Z(n5136) );
  AND U5227 ( .A(n12128), .B(n159), .Z(n5177) );
  XOR U5228 ( .A(n5392), .B(n5393), .Z(n5133) );
  ANDN U5229 ( .A(n5394), .B(n5395), .Z(n5393) );
  XNOR U5230 ( .A(n5392), .B(n5396), .Z(n5394) );
  XOR U5231 ( .A(n5144), .B(n5397), .Z(n5137) );
  IV U5232 ( .A(n5143), .Z(n5397) );
  XNOR U5233 ( .A(n5140), .B(n5170), .Z(n5143) );
  AND U5234 ( .A(n12387), .B(n80), .Z(n5170) );
  XOR U5235 ( .A(n5398), .B(n5399), .Z(n5140) );
  ANDN U5236 ( .A(n5400), .B(n5401), .Z(n5399) );
  XNOR U5237 ( .A(n5398), .B(n5402), .Z(n5400) );
  XOR U5238 ( .A(n5149), .B(n5403), .Z(n5144) );
  IV U5239 ( .A(n5148), .Z(n5403) );
  XNOR U5240 ( .A(n5145), .B(n5404), .Z(n5148) );
  AND U5241 ( .A(n42), .B(n12644), .Z(n5404) );
  XOR U5242 ( .A(n5405), .B(n5406), .Z(n5145) );
  ANDN U5243 ( .A(n5407), .B(n5408), .Z(n5406) );
  XNOR U5244 ( .A(n5405), .B(n5409), .Z(n5407) );
  XNOR U5245 ( .A(n5410), .B(n5411), .Z(n5149) );
  ANDN U5246 ( .A(n5412), .B(n5413), .Z(n5411) );
  XNOR U5247 ( .A(n5410), .B(n5414), .Z(n5412) );
  XNOR U5248 ( .A(n5158), .B(n5150), .Z(n5168) );
  XOR U5249 ( .A(n5415), .B(n5416), .Z(n5150) );
  AND U5250 ( .A(n5417), .B(n5418), .Z(n5416) );
  XNOR U5251 ( .A(n5419), .B(n5415), .Z(n5418) );
  XOR U5252 ( .A(n5156), .B(n5420), .Z(n5158) );
  ANDN U5253 ( .A(n12644), .B(n43), .Z(n5420) );
  XOR U5254 ( .A(n5421), .B(n5422), .Z(n5156) );
  AND U5255 ( .A(n5423), .B(n5424), .Z(n5422) );
  XNOR U5256 ( .A(n5421), .B(n5425), .Z(n5424) );
  XOR U5257 ( .A(n5154), .B(n5164), .Z(n5167) );
  XOR U5258 ( .A(n5426), .B(n5427), .Z(n5154) );
  IV U5259 ( .A(n5428), .Z(n5427) );
  XOR U5260 ( .A(n5429), .B(n5430), .Z(n5164) );
  AND U5261 ( .A(n5429), .B(n5431), .Z(n5430) );
  XOR U5262 ( .A(n5432), .B(n5417), .Z(n5431) );
  XOR U5263 ( .A(n5433), .B(n5425), .Z(n5417) );
  XOR U5264 ( .A(n5175), .B(n5434), .Z(n5425) );
  IV U5265 ( .A(n5174), .Z(n5434) );
  XNOR U5266 ( .A(n5171), .B(n5435), .Z(n5174) );
  XOR U5267 ( .A(n5436), .B(n5437), .Z(n5171) );
  ANDN U5268 ( .A(n5438), .B(n5439), .Z(n5437) );
  XNOR U5269 ( .A(n5436), .B(n5440), .Z(n5438) );
  XOR U5270 ( .A(n5182), .B(n5441), .Z(n5175) );
  IV U5271 ( .A(n5181), .Z(n5441) );
  XNOR U5272 ( .A(n5178), .B(n5442), .Z(n5181) );
  XOR U5273 ( .A(n5443), .B(n5444), .Z(n5178) );
  ANDN U5274 ( .A(n5445), .B(n5446), .Z(n5444) );
  XNOR U5275 ( .A(n5443), .B(n5447), .Z(n5445) );
  XOR U5276 ( .A(n5189), .B(n5448), .Z(n5182) );
  IV U5277 ( .A(n5188), .Z(n5448) );
  XNOR U5278 ( .A(n5185), .B(n5449), .Z(n5188) );
  XOR U5279 ( .A(n5450), .B(n5451), .Z(n5185) );
  ANDN U5280 ( .A(n5452), .B(n5453), .Z(n5451) );
  XNOR U5281 ( .A(n5450), .B(n5454), .Z(n5452) );
  XOR U5282 ( .A(n5196), .B(n5455), .Z(n5189) );
  IV U5283 ( .A(n5195), .Z(n5455) );
  XNOR U5284 ( .A(n5192), .B(n5456), .Z(n5195) );
  XOR U5285 ( .A(n5457), .B(n5458), .Z(n5192) );
  ANDN U5286 ( .A(n5459), .B(n5460), .Z(n5458) );
  XNOR U5287 ( .A(n5457), .B(n5461), .Z(n5459) );
  XOR U5288 ( .A(n5203), .B(n5462), .Z(n5196) );
  IV U5289 ( .A(n5202), .Z(n5462) );
  XNOR U5290 ( .A(n5199), .B(n5463), .Z(n5202) );
  XOR U5291 ( .A(n5464), .B(n5465), .Z(n5199) );
  ANDN U5292 ( .A(n5466), .B(n5467), .Z(n5465) );
  XNOR U5293 ( .A(n5464), .B(n5468), .Z(n5466) );
  XOR U5294 ( .A(n5210), .B(n5469), .Z(n5203) );
  IV U5295 ( .A(n5209), .Z(n5469) );
  XNOR U5296 ( .A(n5206), .B(n5470), .Z(n5209) );
  XOR U5297 ( .A(n5471), .B(n5472), .Z(n5206) );
  ANDN U5298 ( .A(n5473), .B(n5474), .Z(n5472) );
  XNOR U5299 ( .A(n5471), .B(n5475), .Z(n5473) );
  XOR U5300 ( .A(n5217), .B(n5476), .Z(n5210) );
  IV U5301 ( .A(n5216), .Z(n5476) );
  XNOR U5302 ( .A(n5213), .B(n5477), .Z(n5216) );
  XOR U5303 ( .A(n5478), .B(n5479), .Z(n5213) );
  ANDN U5304 ( .A(n5480), .B(n5481), .Z(n5479) );
  XNOR U5305 ( .A(n5478), .B(n5482), .Z(n5480) );
  XOR U5306 ( .A(n5224), .B(n5483), .Z(n5217) );
  IV U5307 ( .A(n5223), .Z(n5483) );
  XNOR U5308 ( .A(n5220), .B(n5484), .Z(n5223) );
  XOR U5309 ( .A(n5485), .B(n5486), .Z(n5220) );
  ANDN U5310 ( .A(n5487), .B(n5488), .Z(n5486) );
  XNOR U5311 ( .A(n5485), .B(n5489), .Z(n5487) );
  XOR U5312 ( .A(n5231), .B(n5490), .Z(n5224) );
  IV U5313 ( .A(n5230), .Z(n5490) );
  XNOR U5314 ( .A(n5227), .B(n5491), .Z(n5230) );
  XOR U5315 ( .A(n5492), .B(n5493), .Z(n5227) );
  ANDN U5316 ( .A(n5494), .B(n5495), .Z(n5493) );
  XNOR U5317 ( .A(n5492), .B(n5496), .Z(n5494) );
  XOR U5318 ( .A(n5238), .B(n5497), .Z(n5231) );
  IV U5319 ( .A(n5237), .Z(n5497) );
  XNOR U5320 ( .A(n5234), .B(n5498), .Z(n5237) );
  XOR U5321 ( .A(n5499), .B(n5500), .Z(n5234) );
  ANDN U5322 ( .A(n5501), .B(n5502), .Z(n5500) );
  XNOR U5323 ( .A(n5499), .B(n5503), .Z(n5501) );
  XOR U5324 ( .A(n5245), .B(n5504), .Z(n5238) );
  IV U5325 ( .A(n5244), .Z(n5504) );
  XNOR U5326 ( .A(n5241), .B(n5505), .Z(n5244) );
  XOR U5327 ( .A(n5506), .B(n5507), .Z(n5241) );
  ANDN U5328 ( .A(n5508), .B(n5509), .Z(n5507) );
  XNOR U5329 ( .A(n5506), .B(n5510), .Z(n5508) );
  XOR U5330 ( .A(n5252), .B(n5511), .Z(n5245) );
  IV U5331 ( .A(n5251), .Z(n5511) );
  XNOR U5332 ( .A(n5248), .B(n5512), .Z(n5251) );
  XOR U5333 ( .A(n5513), .B(n5514), .Z(n5248) );
  ANDN U5334 ( .A(n5515), .B(n5516), .Z(n5514) );
  XNOR U5335 ( .A(n5513), .B(n5517), .Z(n5515) );
  XOR U5336 ( .A(n5259), .B(n5518), .Z(n5252) );
  IV U5337 ( .A(n5258), .Z(n5518) );
  XNOR U5338 ( .A(n5255), .B(n5519), .Z(n5258) );
  XOR U5339 ( .A(n5520), .B(n5521), .Z(n5255) );
  ANDN U5340 ( .A(n5522), .B(n5523), .Z(n5521) );
  XNOR U5341 ( .A(n5520), .B(n5524), .Z(n5522) );
  XOR U5342 ( .A(n5266), .B(n5525), .Z(n5259) );
  IV U5343 ( .A(n5265), .Z(n5525) );
  XNOR U5344 ( .A(n5262), .B(n5526), .Z(n5265) );
  XOR U5345 ( .A(n5527), .B(n5528), .Z(n5262) );
  ANDN U5346 ( .A(n5529), .B(n5530), .Z(n5528) );
  XNOR U5347 ( .A(n5527), .B(n5531), .Z(n5529) );
  XOR U5348 ( .A(n5273), .B(n5532), .Z(n5266) );
  IV U5349 ( .A(n5272), .Z(n5532) );
  XNOR U5350 ( .A(n5269), .B(n5533), .Z(n5272) );
  XOR U5351 ( .A(n5534), .B(n5535), .Z(n5269) );
  ANDN U5352 ( .A(n5536), .B(n5537), .Z(n5535) );
  XNOR U5353 ( .A(n5534), .B(n5538), .Z(n5536) );
  XOR U5354 ( .A(n5280), .B(n5539), .Z(n5273) );
  IV U5355 ( .A(n5279), .Z(n5539) );
  XNOR U5356 ( .A(n5276), .B(n5540), .Z(n5279) );
  XOR U5357 ( .A(n5541), .B(n5542), .Z(n5276) );
  ANDN U5358 ( .A(n5543), .B(n5544), .Z(n5542) );
  XNOR U5359 ( .A(n5541), .B(n5545), .Z(n5543) );
  XOR U5360 ( .A(n5287), .B(n5546), .Z(n5280) );
  IV U5361 ( .A(n5286), .Z(n5546) );
  XNOR U5362 ( .A(n5283), .B(n5547), .Z(n5286) );
  XOR U5363 ( .A(n5548), .B(n5549), .Z(n5283) );
  ANDN U5364 ( .A(n5550), .B(n5551), .Z(n5549) );
  XNOR U5365 ( .A(n5548), .B(n5552), .Z(n5550) );
  XOR U5366 ( .A(n5294), .B(n5553), .Z(n5287) );
  IV U5367 ( .A(n5293), .Z(n5553) );
  XNOR U5368 ( .A(n5290), .B(n5554), .Z(n5293) );
  XOR U5369 ( .A(n5555), .B(n5556), .Z(n5290) );
  ANDN U5370 ( .A(n5557), .B(n5558), .Z(n5556) );
  XNOR U5371 ( .A(n5555), .B(n5559), .Z(n5557) );
  XOR U5372 ( .A(n5300), .B(n5560), .Z(n5294) );
  IV U5373 ( .A(n5299), .Z(n5560) );
  XNOR U5374 ( .A(n5296), .B(n5561), .Z(n5299) );
  XOR U5375 ( .A(n5562), .B(n5563), .Z(n5296) );
  ANDN U5376 ( .A(n5564), .B(n5565), .Z(n5563) );
  XNOR U5377 ( .A(n5562), .B(n5566), .Z(n5564) );
  XOR U5378 ( .A(n5306), .B(n5567), .Z(n5300) );
  IV U5379 ( .A(n5305), .Z(n5567) );
  XNOR U5380 ( .A(n5302), .B(n5554), .Z(n5305) );
  AND U5381 ( .A(n6118), .B(n5030), .Z(n5554) );
  XOR U5382 ( .A(n5568), .B(n5569), .Z(n5302) );
  ANDN U5383 ( .A(n5570), .B(n5571), .Z(n5569) );
  XNOR U5384 ( .A(n5568), .B(n5572), .Z(n5570) );
  XOR U5385 ( .A(n5312), .B(n5573), .Z(n5306) );
  IV U5386 ( .A(n5311), .Z(n5573) );
  XNOR U5387 ( .A(n5308), .B(n5547), .Z(n5311) );
  AND U5388 ( .A(n6688), .B(n4525), .Z(n5547) );
  XOR U5389 ( .A(n5574), .B(n5575), .Z(n5308) );
  ANDN U5390 ( .A(n5576), .B(n5577), .Z(n5575) );
  XNOR U5391 ( .A(n5574), .B(n5578), .Z(n5576) );
  XOR U5392 ( .A(n5318), .B(n5579), .Z(n5312) );
  IV U5393 ( .A(n5317), .Z(n5579) );
  XNOR U5394 ( .A(n5314), .B(n5540), .Z(n5317) );
  AND U5395 ( .A(n7241), .B(n4046), .Z(n5540) );
  XOR U5396 ( .A(n5580), .B(n5581), .Z(n5314) );
  ANDN U5397 ( .A(n5582), .B(n5583), .Z(n5581) );
  XNOR U5398 ( .A(n5580), .B(n5584), .Z(n5582) );
  XOR U5399 ( .A(n5324), .B(n5585), .Z(n5318) );
  IV U5400 ( .A(n5323), .Z(n5585) );
  XNOR U5401 ( .A(n5320), .B(n5533), .Z(n5323) );
  AND U5402 ( .A(n7770), .B(n3593), .Z(n5533) );
  XOR U5403 ( .A(n5586), .B(n5587), .Z(n5320) );
  ANDN U5404 ( .A(n5588), .B(n5589), .Z(n5587) );
  XNOR U5405 ( .A(n5586), .B(n5590), .Z(n5588) );
  XOR U5406 ( .A(n5330), .B(n5591), .Z(n5324) );
  IV U5407 ( .A(n5329), .Z(n5591) );
  XNOR U5408 ( .A(n5326), .B(n5526), .Z(n5329) );
  AND U5409 ( .A(n8272), .B(n3166), .Z(n5526) );
  XOR U5410 ( .A(n5592), .B(n5593), .Z(n5326) );
  ANDN U5411 ( .A(n5594), .B(n5595), .Z(n5593) );
  XNOR U5412 ( .A(n5592), .B(n5596), .Z(n5594) );
  XOR U5413 ( .A(n5336), .B(n5597), .Z(n5330) );
  IV U5414 ( .A(n5335), .Z(n5597) );
  XNOR U5415 ( .A(n5332), .B(n5519), .Z(n5335) );
  AND U5416 ( .A(n8748), .B(n2765), .Z(n5519) );
  XOR U5417 ( .A(n5598), .B(n5599), .Z(n5332) );
  ANDN U5418 ( .A(n5600), .B(n5601), .Z(n5599) );
  XNOR U5419 ( .A(n5598), .B(n5602), .Z(n5600) );
  XOR U5420 ( .A(n5342), .B(n5603), .Z(n5336) );
  IV U5421 ( .A(n5341), .Z(n5603) );
  XNOR U5422 ( .A(n5338), .B(n5512), .Z(n5341) );
  AND U5423 ( .A(n9198), .B(n2396), .Z(n5512) );
  XOR U5424 ( .A(n5604), .B(n5605), .Z(n5338) );
  ANDN U5425 ( .A(n5606), .B(n5607), .Z(n5605) );
  XNOR U5426 ( .A(n5604), .B(n5608), .Z(n5606) );
  XOR U5427 ( .A(n5348), .B(n5609), .Z(n5342) );
  IV U5428 ( .A(n5347), .Z(n5609) );
  XNOR U5429 ( .A(n5344), .B(n5505), .Z(n5347) );
  AND U5430 ( .A(n9621), .B(n2053), .Z(n5505) );
  XOR U5431 ( .A(n5610), .B(n5611), .Z(n5344) );
  ANDN U5432 ( .A(n5612), .B(n5613), .Z(n5611) );
  XNOR U5433 ( .A(n5610), .B(n5614), .Z(n5612) );
  XOR U5434 ( .A(n5354), .B(n5615), .Z(n5348) );
  IV U5435 ( .A(n5353), .Z(n5615) );
  XNOR U5436 ( .A(n5350), .B(n5498), .Z(n5353) );
  AND U5437 ( .A(n10017), .B(n1737), .Z(n5498) );
  XOR U5438 ( .A(n5616), .B(n5617), .Z(n5350) );
  ANDN U5439 ( .A(n5618), .B(n5619), .Z(n5617) );
  XNOR U5440 ( .A(n5616), .B(n5620), .Z(n5618) );
  XOR U5441 ( .A(n5360), .B(n5621), .Z(n5354) );
  IV U5442 ( .A(n5359), .Z(n5621) );
  XNOR U5443 ( .A(n5356), .B(n5491), .Z(n5359) );
  AND U5444 ( .A(n10387), .B(n1448), .Z(n5491) );
  XOR U5445 ( .A(n5622), .B(n5623), .Z(n5356) );
  ANDN U5446 ( .A(n5624), .B(n5625), .Z(n5623) );
  XNOR U5447 ( .A(n5622), .B(n5626), .Z(n5624) );
  XOR U5448 ( .A(n5366), .B(n5627), .Z(n5360) );
  IV U5449 ( .A(n5365), .Z(n5627) );
  XNOR U5450 ( .A(n5362), .B(n5484), .Z(n5365) );
  AND U5451 ( .A(n10731), .B(n1185), .Z(n5484) );
  XOR U5452 ( .A(n5628), .B(n5629), .Z(n5362) );
  ANDN U5453 ( .A(n5630), .B(n5631), .Z(n5629) );
  XNOR U5454 ( .A(n5628), .B(n5632), .Z(n5630) );
  XOR U5455 ( .A(n5372), .B(n5633), .Z(n5366) );
  IV U5456 ( .A(n5371), .Z(n5633) );
  XNOR U5457 ( .A(n5368), .B(n5477), .Z(n5371) );
  AND U5458 ( .A(n11049), .B(n948), .Z(n5477) );
  XOR U5459 ( .A(n5634), .B(n5635), .Z(n5368) );
  ANDN U5460 ( .A(n5636), .B(n5637), .Z(n5635) );
  XNOR U5461 ( .A(n5634), .B(n5638), .Z(n5636) );
  XOR U5462 ( .A(n5378), .B(n5639), .Z(n5372) );
  IV U5463 ( .A(n5377), .Z(n5639) );
  XNOR U5464 ( .A(n5374), .B(n5470), .Z(n5377) );
  AND U5465 ( .A(n11341), .B(n736), .Z(n5470) );
  XOR U5466 ( .A(n5640), .B(n5641), .Z(n5374) );
  ANDN U5467 ( .A(n5642), .B(n5643), .Z(n5641) );
  XNOR U5468 ( .A(n5640), .B(n5644), .Z(n5642) );
  XOR U5469 ( .A(n5384), .B(n5645), .Z(n5378) );
  IV U5470 ( .A(n5383), .Z(n5645) );
  XNOR U5471 ( .A(n5380), .B(n5463), .Z(n5383) );
  AND U5472 ( .A(n11607), .B(n552), .Z(n5463) );
  XOR U5473 ( .A(n5646), .B(n5647), .Z(n5380) );
  ANDN U5474 ( .A(n5648), .B(n5649), .Z(n5647) );
  XNOR U5475 ( .A(n5646), .B(n5650), .Z(n5648) );
  XOR U5476 ( .A(n5390), .B(n5651), .Z(n5384) );
  IV U5477 ( .A(n5389), .Z(n5651) );
  XNOR U5478 ( .A(n5386), .B(n5456), .Z(n5389) );
  AND U5479 ( .A(n11869), .B(n395), .Z(n5456) );
  XOR U5480 ( .A(n5652), .B(n5653), .Z(n5386) );
  ANDN U5481 ( .A(n5654), .B(n5655), .Z(n5653) );
  XNOR U5482 ( .A(n5652), .B(n5656), .Z(n5654) );
  XOR U5483 ( .A(n5396), .B(n5657), .Z(n5390) );
  IV U5484 ( .A(n5395), .Z(n5657) );
  XNOR U5485 ( .A(n5392), .B(n5449), .Z(n5395) );
  AND U5486 ( .A(n12128), .B(n264), .Z(n5449) );
  XOR U5487 ( .A(n5658), .B(n5659), .Z(n5392) );
  ANDN U5488 ( .A(n5660), .B(n5661), .Z(n5659) );
  XNOR U5489 ( .A(n5658), .B(n5662), .Z(n5660) );
  XOR U5490 ( .A(n5402), .B(n5663), .Z(n5396) );
  IV U5491 ( .A(n5401), .Z(n5663) );
  XNOR U5492 ( .A(n5398), .B(n5442), .Z(n5401) );
  AND U5493 ( .A(n12387), .B(n159), .Z(n5442) );
  XOR U5494 ( .A(n5664), .B(n5665), .Z(n5398) );
  ANDN U5495 ( .A(n5666), .B(n5667), .Z(n5665) );
  XNOR U5496 ( .A(n5664), .B(n5668), .Z(n5666) );
  XOR U5497 ( .A(n5409), .B(n5669), .Z(n5402) );
  IV U5498 ( .A(n5408), .Z(n5669) );
  XNOR U5499 ( .A(n5405), .B(n5435), .Z(n5408) );
  AND U5500 ( .A(n12644), .B(n80), .Z(n5435) );
  XOR U5501 ( .A(n5670), .B(n5671), .Z(n5405) );
  ANDN U5502 ( .A(n5672), .B(n5673), .Z(n5671) );
  XNOR U5503 ( .A(n5670), .B(n5674), .Z(n5672) );
  XOR U5504 ( .A(n5414), .B(n5675), .Z(n5409) );
  IV U5505 ( .A(n5413), .Z(n5675) );
  XNOR U5506 ( .A(n5410), .B(n5676), .Z(n5413) );
  AND U5507 ( .A(n42), .B(n12880), .Z(n5676) );
  XOR U5508 ( .A(n5677), .B(n5678), .Z(n5410) );
  ANDN U5509 ( .A(n5679), .B(n5680), .Z(n5678) );
  XNOR U5510 ( .A(n5677), .B(n5681), .Z(n5679) );
  XNOR U5511 ( .A(n5682), .B(n5683), .Z(n5414) );
  ANDN U5512 ( .A(n5684), .B(n5685), .Z(n5683) );
  XNOR U5513 ( .A(n5682), .B(n5686), .Z(n5684) );
  XNOR U5514 ( .A(n5423), .B(n5415), .Z(n5433) );
  XOR U5515 ( .A(n5687), .B(n5688), .Z(n5415) );
  AND U5516 ( .A(n5689), .B(n5690), .Z(n5688) );
  XNOR U5517 ( .A(n5691), .B(n5687), .Z(n5690) );
  XOR U5518 ( .A(n5421), .B(n5692), .Z(n5423) );
  ANDN U5519 ( .A(n12880), .B(n43), .Z(n5692) );
  XOR U5520 ( .A(n5693), .B(n5694), .Z(n5421) );
  AND U5521 ( .A(n5695), .B(n5696), .Z(n5694) );
  XNOR U5522 ( .A(n5693), .B(n5697), .Z(n5696) );
  XOR U5523 ( .A(n5419), .B(n5429), .Z(n5432) );
  XOR U5524 ( .A(n5698), .B(n5699), .Z(n5419) );
  IV U5525 ( .A(n5700), .Z(n5699) );
  XOR U5526 ( .A(n5701), .B(n5702), .Z(n5429) );
  AND U5527 ( .A(n5701), .B(n5703), .Z(n5702) );
  XOR U5528 ( .A(n5704), .B(n5689), .Z(n5703) );
  XOR U5529 ( .A(n5705), .B(n5697), .Z(n5689) );
  XOR U5530 ( .A(n5440), .B(n5706), .Z(n5697) );
  IV U5531 ( .A(n5439), .Z(n5706) );
  XNOR U5532 ( .A(n5436), .B(n5707), .Z(n5439) );
  XOR U5533 ( .A(n5708), .B(n5709), .Z(n5436) );
  ANDN U5534 ( .A(n5710), .B(n5711), .Z(n5709) );
  XNOR U5535 ( .A(n5708), .B(n5712), .Z(n5710) );
  XOR U5536 ( .A(n5447), .B(n5713), .Z(n5440) );
  IV U5537 ( .A(n5446), .Z(n5713) );
  XNOR U5538 ( .A(n5443), .B(n5714), .Z(n5446) );
  XOR U5539 ( .A(n5715), .B(n5716), .Z(n5443) );
  ANDN U5540 ( .A(n5717), .B(n5718), .Z(n5716) );
  XNOR U5541 ( .A(n5715), .B(n5719), .Z(n5717) );
  XOR U5542 ( .A(n5454), .B(n5720), .Z(n5447) );
  IV U5543 ( .A(n5453), .Z(n5720) );
  XNOR U5544 ( .A(n5450), .B(n5721), .Z(n5453) );
  XOR U5545 ( .A(n5722), .B(n5723), .Z(n5450) );
  ANDN U5546 ( .A(n5724), .B(n5725), .Z(n5723) );
  XNOR U5547 ( .A(n5722), .B(n5726), .Z(n5724) );
  XOR U5548 ( .A(n5461), .B(n5727), .Z(n5454) );
  IV U5549 ( .A(n5460), .Z(n5727) );
  XNOR U5550 ( .A(n5457), .B(n5728), .Z(n5460) );
  XOR U5551 ( .A(n5729), .B(n5730), .Z(n5457) );
  ANDN U5552 ( .A(n5731), .B(n5732), .Z(n5730) );
  XNOR U5553 ( .A(n5729), .B(n5733), .Z(n5731) );
  XOR U5554 ( .A(n5468), .B(n5734), .Z(n5461) );
  IV U5555 ( .A(n5467), .Z(n5734) );
  XNOR U5556 ( .A(n5464), .B(n5735), .Z(n5467) );
  XOR U5557 ( .A(n5736), .B(n5737), .Z(n5464) );
  ANDN U5558 ( .A(n5738), .B(n5739), .Z(n5737) );
  XNOR U5559 ( .A(n5736), .B(n5740), .Z(n5738) );
  XOR U5560 ( .A(n5475), .B(n5741), .Z(n5468) );
  IV U5561 ( .A(n5474), .Z(n5741) );
  XNOR U5562 ( .A(n5471), .B(n5742), .Z(n5474) );
  XOR U5563 ( .A(n5743), .B(n5744), .Z(n5471) );
  ANDN U5564 ( .A(n5745), .B(n5746), .Z(n5744) );
  XNOR U5565 ( .A(n5743), .B(n5747), .Z(n5745) );
  XOR U5566 ( .A(n5482), .B(n5748), .Z(n5475) );
  IV U5567 ( .A(n5481), .Z(n5748) );
  XNOR U5568 ( .A(n5478), .B(n5749), .Z(n5481) );
  XOR U5569 ( .A(n5750), .B(n5751), .Z(n5478) );
  ANDN U5570 ( .A(n5752), .B(n5753), .Z(n5751) );
  XNOR U5571 ( .A(n5750), .B(n5754), .Z(n5752) );
  XOR U5572 ( .A(n5489), .B(n5755), .Z(n5482) );
  IV U5573 ( .A(n5488), .Z(n5755) );
  XNOR U5574 ( .A(n5485), .B(n5756), .Z(n5488) );
  XOR U5575 ( .A(n5757), .B(n5758), .Z(n5485) );
  ANDN U5576 ( .A(n5759), .B(n5760), .Z(n5758) );
  XNOR U5577 ( .A(n5757), .B(n5761), .Z(n5759) );
  XOR U5578 ( .A(n5496), .B(n5762), .Z(n5489) );
  IV U5579 ( .A(n5495), .Z(n5762) );
  XNOR U5580 ( .A(n5492), .B(n5763), .Z(n5495) );
  XOR U5581 ( .A(n5764), .B(n5765), .Z(n5492) );
  ANDN U5582 ( .A(n5766), .B(n5767), .Z(n5765) );
  XNOR U5583 ( .A(n5764), .B(n5768), .Z(n5766) );
  XOR U5584 ( .A(n5503), .B(n5769), .Z(n5496) );
  IV U5585 ( .A(n5502), .Z(n5769) );
  XNOR U5586 ( .A(n5499), .B(n5770), .Z(n5502) );
  XOR U5587 ( .A(n5771), .B(n5772), .Z(n5499) );
  ANDN U5588 ( .A(n5773), .B(n5774), .Z(n5772) );
  XNOR U5589 ( .A(n5771), .B(n5775), .Z(n5773) );
  XOR U5590 ( .A(n5510), .B(n5776), .Z(n5503) );
  IV U5591 ( .A(n5509), .Z(n5776) );
  XNOR U5592 ( .A(n5506), .B(n5777), .Z(n5509) );
  XOR U5593 ( .A(n5778), .B(n5779), .Z(n5506) );
  ANDN U5594 ( .A(n5780), .B(n5781), .Z(n5779) );
  XNOR U5595 ( .A(n5778), .B(n5782), .Z(n5780) );
  XOR U5596 ( .A(n5517), .B(n5783), .Z(n5510) );
  IV U5597 ( .A(n5516), .Z(n5783) );
  XNOR U5598 ( .A(n5513), .B(n5784), .Z(n5516) );
  XOR U5599 ( .A(n5785), .B(n5786), .Z(n5513) );
  ANDN U5600 ( .A(n5787), .B(n5788), .Z(n5786) );
  XNOR U5601 ( .A(n5785), .B(n5789), .Z(n5787) );
  XOR U5602 ( .A(n5524), .B(n5790), .Z(n5517) );
  IV U5603 ( .A(n5523), .Z(n5790) );
  XNOR U5604 ( .A(n5520), .B(n5791), .Z(n5523) );
  XOR U5605 ( .A(n5792), .B(n5793), .Z(n5520) );
  ANDN U5606 ( .A(n5794), .B(n5795), .Z(n5793) );
  XNOR U5607 ( .A(n5792), .B(n5796), .Z(n5794) );
  XOR U5608 ( .A(n5531), .B(n5797), .Z(n5524) );
  IV U5609 ( .A(n5530), .Z(n5797) );
  XNOR U5610 ( .A(n5527), .B(n5798), .Z(n5530) );
  XOR U5611 ( .A(n5799), .B(n5800), .Z(n5527) );
  ANDN U5612 ( .A(n5801), .B(n5802), .Z(n5800) );
  XNOR U5613 ( .A(n5799), .B(n5803), .Z(n5801) );
  XOR U5614 ( .A(n5538), .B(n5804), .Z(n5531) );
  IV U5615 ( .A(n5537), .Z(n5804) );
  XNOR U5616 ( .A(n5534), .B(n5805), .Z(n5537) );
  XOR U5617 ( .A(n5806), .B(n5807), .Z(n5534) );
  ANDN U5618 ( .A(n5808), .B(n5809), .Z(n5807) );
  XNOR U5619 ( .A(n5806), .B(n5810), .Z(n5808) );
  XOR U5620 ( .A(n5545), .B(n5811), .Z(n5538) );
  IV U5621 ( .A(n5544), .Z(n5811) );
  XNOR U5622 ( .A(n5541), .B(n5812), .Z(n5544) );
  XOR U5623 ( .A(n5813), .B(n5814), .Z(n5541) );
  ANDN U5624 ( .A(n5815), .B(n5816), .Z(n5814) );
  XNOR U5625 ( .A(n5813), .B(n5817), .Z(n5815) );
  XOR U5626 ( .A(n5552), .B(n5818), .Z(n5545) );
  IV U5627 ( .A(n5551), .Z(n5818) );
  XNOR U5628 ( .A(n5548), .B(n5819), .Z(n5551) );
  XOR U5629 ( .A(n5820), .B(n5821), .Z(n5548) );
  ANDN U5630 ( .A(n5822), .B(n5823), .Z(n5821) );
  XNOR U5631 ( .A(n5820), .B(n5824), .Z(n5822) );
  XOR U5632 ( .A(n5559), .B(n5825), .Z(n5552) );
  IV U5633 ( .A(n5558), .Z(n5825) );
  XNOR U5634 ( .A(n5555), .B(n5826), .Z(n5558) );
  XOR U5635 ( .A(n5827), .B(n5828), .Z(n5555) );
  ANDN U5636 ( .A(n5829), .B(n5830), .Z(n5828) );
  XNOR U5637 ( .A(n5827), .B(n5831), .Z(n5829) );
  XOR U5638 ( .A(n5566), .B(n5832), .Z(n5559) );
  IV U5639 ( .A(n5565), .Z(n5832) );
  XNOR U5640 ( .A(n5562), .B(n5833), .Z(n5565) );
  XOR U5641 ( .A(n5834), .B(n5835), .Z(n5562) );
  ANDN U5642 ( .A(n5836), .B(n5837), .Z(n5835) );
  XNOR U5643 ( .A(n5834), .B(n5838), .Z(n5836) );
  XOR U5644 ( .A(n5572), .B(n5839), .Z(n5566) );
  IV U5645 ( .A(n5571), .Z(n5839) );
  XNOR U5646 ( .A(n5568), .B(n5833), .Z(n5571) );
  AND U5647 ( .A(n6118), .B(n5561), .Z(n5833) );
  XOR U5648 ( .A(n5840), .B(n5841), .Z(n5568) );
  ANDN U5649 ( .A(n5842), .B(n5843), .Z(n5841) );
  XNOR U5650 ( .A(n5840), .B(n5844), .Z(n5842) );
  XOR U5651 ( .A(n5578), .B(n5845), .Z(n5572) );
  IV U5652 ( .A(n5577), .Z(n5845) );
  XNOR U5653 ( .A(n5574), .B(n5826), .Z(n5577) );
  AND U5654 ( .A(n6688), .B(n5030), .Z(n5826) );
  XOR U5655 ( .A(n5846), .B(n5847), .Z(n5574) );
  ANDN U5656 ( .A(n5848), .B(n5849), .Z(n5847) );
  XNOR U5657 ( .A(n5846), .B(n5850), .Z(n5848) );
  XOR U5658 ( .A(n5584), .B(n5851), .Z(n5578) );
  IV U5659 ( .A(n5583), .Z(n5851) );
  XNOR U5660 ( .A(n5580), .B(n5819), .Z(n5583) );
  AND U5661 ( .A(n7241), .B(n4525), .Z(n5819) );
  XOR U5662 ( .A(n5852), .B(n5853), .Z(n5580) );
  ANDN U5663 ( .A(n5854), .B(n5855), .Z(n5853) );
  XNOR U5664 ( .A(n5852), .B(n5856), .Z(n5854) );
  XOR U5665 ( .A(n5590), .B(n5857), .Z(n5584) );
  IV U5666 ( .A(n5589), .Z(n5857) );
  XNOR U5667 ( .A(n5586), .B(n5812), .Z(n5589) );
  AND U5668 ( .A(n7770), .B(n4046), .Z(n5812) );
  XOR U5669 ( .A(n5858), .B(n5859), .Z(n5586) );
  ANDN U5670 ( .A(n5860), .B(n5861), .Z(n5859) );
  XNOR U5671 ( .A(n5858), .B(n5862), .Z(n5860) );
  XOR U5672 ( .A(n5596), .B(n5863), .Z(n5590) );
  IV U5673 ( .A(n5595), .Z(n5863) );
  XNOR U5674 ( .A(n5592), .B(n5805), .Z(n5595) );
  AND U5675 ( .A(n8272), .B(n3593), .Z(n5805) );
  XOR U5676 ( .A(n5864), .B(n5865), .Z(n5592) );
  ANDN U5677 ( .A(n5866), .B(n5867), .Z(n5865) );
  XNOR U5678 ( .A(n5864), .B(n5868), .Z(n5866) );
  XOR U5679 ( .A(n5602), .B(n5869), .Z(n5596) );
  IV U5680 ( .A(n5601), .Z(n5869) );
  XNOR U5681 ( .A(n5598), .B(n5798), .Z(n5601) );
  AND U5682 ( .A(n8748), .B(n3166), .Z(n5798) );
  XOR U5683 ( .A(n5870), .B(n5871), .Z(n5598) );
  ANDN U5684 ( .A(n5872), .B(n5873), .Z(n5871) );
  XNOR U5685 ( .A(n5870), .B(n5874), .Z(n5872) );
  XOR U5686 ( .A(n5608), .B(n5875), .Z(n5602) );
  IV U5687 ( .A(n5607), .Z(n5875) );
  XNOR U5688 ( .A(n5604), .B(n5791), .Z(n5607) );
  AND U5689 ( .A(n9198), .B(n2765), .Z(n5791) );
  XOR U5690 ( .A(n5876), .B(n5877), .Z(n5604) );
  ANDN U5691 ( .A(n5878), .B(n5879), .Z(n5877) );
  XNOR U5692 ( .A(n5876), .B(n5880), .Z(n5878) );
  XOR U5693 ( .A(n5614), .B(n5881), .Z(n5608) );
  IV U5694 ( .A(n5613), .Z(n5881) );
  XNOR U5695 ( .A(n5610), .B(n5784), .Z(n5613) );
  AND U5696 ( .A(n9621), .B(n2396), .Z(n5784) );
  XOR U5697 ( .A(n5882), .B(n5883), .Z(n5610) );
  ANDN U5698 ( .A(n5884), .B(n5885), .Z(n5883) );
  XNOR U5699 ( .A(n5882), .B(n5886), .Z(n5884) );
  XOR U5700 ( .A(n5620), .B(n5887), .Z(n5614) );
  IV U5701 ( .A(n5619), .Z(n5887) );
  XNOR U5702 ( .A(n5616), .B(n5777), .Z(n5619) );
  AND U5703 ( .A(n10017), .B(n2053), .Z(n5777) );
  XOR U5704 ( .A(n5888), .B(n5889), .Z(n5616) );
  ANDN U5705 ( .A(n5890), .B(n5891), .Z(n5889) );
  XNOR U5706 ( .A(n5888), .B(n5892), .Z(n5890) );
  XOR U5707 ( .A(n5626), .B(n5893), .Z(n5620) );
  IV U5708 ( .A(n5625), .Z(n5893) );
  XNOR U5709 ( .A(n5622), .B(n5770), .Z(n5625) );
  AND U5710 ( .A(n10387), .B(n1737), .Z(n5770) );
  XOR U5711 ( .A(n5894), .B(n5895), .Z(n5622) );
  ANDN U5712 ( .A(n5896), .B(n5897), .Z(n5895) );
  XNOR U5713 ( .A(n5894), .B(n5898), .Z(n5896) );
  XOR U5714 ( .A(n5632), .B(n5899), .Z(n5626) );
  IV U5715 ( .A(n5631), .Z(n5899) );
  XNOR U5716 ( .A(n5628), .B(n5763), .Z(n5631) );
  AND U5717 ( .A(n10731), .B(n1448), .Z(n5763) );
  XOR U5718 ( .A(n5900), .B(n5901), .Z(n5628) );
  ANDN U5719 ( .A(n5902), .B(n5903), .Z(n5901) );
  XNOR U5720 ( .A(n5900), .B(n5904), .Z(n5902) );
  XOR U5721 ( .A(n5638), .B(n5905), .Z(n5632) );
  IV U5722 ( .A(n5637), .Z(n5905) );
  XNOR U5723 ( .A(n5634), .B(n5756), .Z(n5637) );
  AND U5724 ( .A(n11049), .B(n1185), .Z(n5756) );
  XOR U5725 ( .A(n5906), .B(n5907), .Z(n5634) );
  ANDN U5726 ( .A(n5908), .B(n5909), .Z(n5907) );
  XNOR U5727 ( .A(n5906), .B(n5910), .Z(n5908) );
  XOR U5728 ( .A(n5644), .B(n5911), .Z(n5638) );
  IV U5729 ( .A(n5643), .Z(n5911) );
  XNOR U5730 ( .A(n5640), .B(n5749), .Z(n5643) );
  AND U5731 ( .A(n11341), .B(n948), .Z(n5749) );
  XOR U5732 ( .A(n5912), .B(n5913), .Z(n5640) );
  ANDN U5733 ( .A(n5914), .B(n5915), .Z(n5913) );
  XNOR U5734 ( .A(n5912), .B(n5916), .Z(n5914) );
  XOR U5735 ( .A(n5650), .B(n5917), .Z(n5644) );
  IV U5736 ( .A(n5649), .Z(n5917) );
  XNOR U5737 ( .A(n5646), .B(n5742), .Z(n5649) );
  AND U5738 ( .A(n11607), .B(n736), .Z(n5742) );
  XOR U5739 ( .A(n5918), .B(n5919), .Z(n5646) );
  ANDN U5740 ( .A(n5920), .B(n5921), .Z(n5919) );
  XNOR U5741 ( .A(n5918), .B(n5922), .Z(n5920) );
  XOR U5742 ( .A(n5656), .B(n5923), .Z(n5650) );
  IV U5743 ( .A(n5655), .Z(n5923) );
  XNOR U5744 ( .A(n5652), .B(n5735), .Z(n5655) );
  AND U5745 ( .A(n11869), .B(n552), .Z(n5735) );
  XOR U5746 ( .A(n5924), .B(n5925), .Z(n5652) );
  ANDN U5747 ( .A(n5926), .B(n5927), .Z(n5925) );
  XNOR U5748 ( .A(n5924), .B(n5928), .Z(n5926) );
  XOR U5749 ( .A(n5662), .B(n5929), .Z(n5656) );
  IV U5750 ( .A(n5661), .Z(n5929) );
  XNOR U5751 ( .A(n5658), .B(n5728), .Z(n5661) );
  AND U5752 ( .A(n12128), .B(n395), .Z(n5728) );
  XOR U5753 ( .A(n5930), .B(n5931), .Z(n5658) );
  ANDN U5754 ( .A(n5932), .B(n5933), .Z(n5931) );
  XNOR U5755 ( .A(n5930), .B(n5934), .Z(n5932) );
  XOR U5756 ( .A(n5668), .B(n5935), .Z(n5662) );
  IV U5757 ( .A(n5667), .Z(n5935) );
  XNOR U5758 ( .A(n5664), .B(n5721), .Z(n5667) );
  AND U5759 ( .A(n12387), .B(n264), .Z(n5721) );
  XOR U5760 ( .A(n5936), .B(n5937), .Z(n5664) );
  ANDN U5761 ( .A(n5938), .B(n5939), .Z(n5937) );
  XNOR U5762 ( .A(n5936), .B(n5940), .Z(n5938) );
  XOR U5763 ( .A(n5674), .B(n5941), .Z(n5668) );
  IV U5764 ( .A(n5673), .Z(n5941) );
  XNOR U5765 ( .A(n5670), .B(n5714), .Z(n5673) );
  AND U5766 ( .A(n12644), .B(n159), .Z(n5714) );
  XOR U5767 ( .A(n5942), .B(n5943), .Z(n5670) );
  ANDN U5768 ( .A(n5944), .B(n5945), .Z(n5943) );
  XNOR U5769 ( .A(n5942), .B(n5946), .Z(n5944) );
  XOR U5770 ( .A(n5681), .B(n5947), .Z(n5674) );
  IV U5771 ( .A(n5680), .Z(n5947) );
  XNOR U5772 ( .A(n5677), .B(n5707), .Z(n5680) );
  AND U5773 ( .A(n12880), .B(n80), .Z(n5707) );
  XOR U5774 ( .A(n5948), .B(n5949), .Z(n5677) );
  ANDN U5775 ( .A(n5950), .B(n5951), .Z(n5949) );
  XNOR U5776 ( .A(n5948), .B(n5952), .Z(n5950) );
  XOR U5777 ( .A(n5686), .B(n5953), .Z(n5681) );
  IV U5778 ( .A(n5685), .Z(n5953) );
  XNOR U5779 ( .A(n5682), .B(n5954), .Z(n5685) );
  AND U5780 ( .A(n42), .B(n13070), .Z(n5954) );
  XOR U5781 ( .A(n5955), .B(n5956), .Z(n5682) );
  ANDN U5782 ( .A(n5957), .B(n5958), .Z(n5956) );
  XNOR U5783 ( .A(n5955), .B(n5959), .Z(n5957) );
  XNOR U5784 ( .A(n5960), .B(n5961), .Z(n5686) );
  ANDN U5785 ( .A(n5962), .B(n5963), .Z(n5961) );
  XNOR U5786 ( .A(n5960), .B(n5964), .Z(n5962) );
  XNOR U5787 ( .A(n5695), .B(n5687), .Z(n5705) );
  XOR U5788 ( .A(n5965), .B(n5966), .Z(n5687) );
  AND U5789 ( .A(n5967), .B(n5968), .Z(n5966) );
  XNOR U5790 ( .A(n5969), .B(n5965), .Z(n5968) );
  XOR U5791 ( .A(n5693), .B(n5970), .Z(n5695) );
  ANDN U5792 ( .A(n13070), .B(n43), .Z(n5970) );
  XOR U5793 ( .A(n5971), .B(n5972), .Z(n5693) );
  AND U5794 ( .A(n5973), .B(n5974), .Z(n5972) );
  XNOR U5795 ( .A(n5971), .B(n5975), .Z(n5974) );
  XOR U5796 ( .A(n5691), .B(n5701), .Z(n5704) );
  XOR U5797 ( .A(n5976), .B(n5977), .Z(n5691) );
  IV U5798 ( .A(n5978), .Z(n5977) );
  XOR U5799 ( .A(n5979), .B(n5980), .Z(n5701) );
  AND U5800 ( .A(n5979), .B(n5981), .Z(n5980) );
  XOR U5801 ( .A(n5982), .B(n5967), .Z(n5981) );
  XOR U5802 ( .A(n5983), .B(n5975), .Z(n5967) );
  XOR U5803 ( .A(n5712), .B(n5984), .Z(n5975) );
  IV U5804 ( .A(n5711), .Z(n5984) );
  XNOR U5805 ( .A(n5708), .B(n5985), .Z(n5711) );
  XOR U5806 ( .A(n5986), .B(n5987), .Z(n5708) );
  ANDN U5807 ( .A(n5988), .B(n5989), .Z(n5987) );
  XNOR U5808 ( .A(n5986), .B(n5990), .Z(n5988) );
  XOR U5809 ( .A(n5719), .B(n5991), .Z(n5712) );
  IV U5810 ( .A(n5718), .Z(n5991) );
  XNOR U5811 ( .A(n5715), .B(n5992), .Z(n5718) );
  XOR U5812 ( .A(n5993), .B(n5994), .Z(n5715) );
  ANDN U5813 ( .A(n5995), .B(n5996), .Z(n5994) );
  XNOR U5814 ( .A(n5993), .B(n5997), .Z(n5995) );
  XOR U5815 ( .A(n5726), .B(n5998), .Z(n5719) );
  IV U5816 ( .A(n5725), .Z(n5998) );
  XNOR U5817 ( .A(n5722), .B(n5999), .Z(n5725) );
  XOR U5818 ( .A(n6000), .B(n6001), .Z(n5722) );
  ANDN U5819 ( .A(n6002), .B(n6003), .Z(n6001) );
  XNOR U5820 ( .A(n6000), .B(n6004), .Z(n6002) );
  XOR U5821 ( .A(n5733), .B(n6005), .Z(n5726) );
  IV U5822 ( .A(n5732), .Z(n6005) );
  XNOR U5823 ( .A(n5729), .B(n6006), .Z(n5732) );
  XOR U5824 ( .A(n6007), .B(n6008), .Z(n5729) );
  ANDN U5825 ( .A(n6009), .B(n6010), .Z(n6008) );
  XNOR U5826 ( .A(n6007), .B(n6011), .Z(n6009) );
  XOR U5827 ( .A(n5740), .B(n6012), .Z(n5733) );
  IV U5828 ( .A(n5739), .Z(n6012) );
  XNOR U5829 ( .A(n5736), .B(n6013), .Z(n5739) );
  XOR U5830 ( .A(n6014), .B(n6015), .Z(n5736) );
  ANDN U5831 ( .A(n6016), .B(n6017), .Z(n6015) );
  XNOR U5832 ( .A(n6014), .B(n6018), .Z(n6016) );
  XOR U5833 ( .A(n5747), .B(n6019), .Z(n5740) );
  IV U5834 ( .A(n5746), .Z(n6019) );
  XNOR U5835 ( .A(n5743), .B(n6020), .Z(n5746) );
  XOR U5836 ( .A(n6021), .B(n6022), .Z(n5743) );
  ANDN U5837 ( .A(n6023), .B(n6024), .Z(n6022) );
  XNOR U5838 ( .A(n6021), .B(n6025), .Z(n6023) );
  XOR U5839 ( .A(n5754), .B(n6026), .Z(n5747) );
  IV U5840 ( .A(n5753), .Z(n6026) );
  XNOR U5841 ( .A(n5750), .B(n6027), .Z(n5753) );
  XOR U5842 ( .A(n6028), .B(n6029), .Z(n5750) );
  ANDN U5843 ( .A(n6030), .B(n6031), .Z(n6029) );
  XNOR U5844 ( .A(n6028), .B(n6032), .Z(n6030) );
  XOR U5845 ( .A(n5761), .B(n6033), .Z(n5754) );
  IV U5846 ( .A(n5760), .Z(n6033) );
  XNOR U5847 ( .A(n5757), .B(n6034), .Z(n5760) );
  XOR U5848 ( .A(n6035), .B(n6036), .Z(n5757) );
  ANDN U5849 ( .A(n6037), .B(n6038), .Z(n6036) );
  XNOR U5850 ( .A(n6035), .B(n6039), .Z(n6037) );
  XOR U5851 ( .A(n5768), .B(n6040), .Z(n5761) );
  IV U5852 ( .A(n5767), .Z(n6040) );
  XNOR U5853 ( .A(n5764), .B(n6041), .Z(n5767) );
  XOR U5854 ( .A(n6042), .B(n6043), .Z(n5764) );
  ANDN U5855 ( .A(n6044), .B(n6045), .Z(n6043) );
  XNOR U5856 ( .A(n6042), .B(n6046), .Z(n6044) );
  XOR U5857 ( .A(n5775), .B(n6047), .Z(n5768) );
  IV U5858 ( .A(n5774), .Z(n6047) );
  XNOR U5859 ( .A(n5771), .B(n6048), .Z(n5774) );
  XOR U5860 ( .A(n6049), .B(n6050), .Z(n5771) );
  ANDN U5861 ( .A(n6051), .B(n6052), .Z(n6050) );
  XNOR U5862 ( .A(n6049), .B(n6053), .Z(n6051) );
  XOR U5863 ( .A(n5782), .B(n6054), .Z(n5775) );
  IV U5864 ( .A(n5781), .Z(n6054) );
  XNOR U5865 ( .A(n5778), .B(n6055), .Z(n5781) );
  XOR U5866 ( .A(n6056), .B(n6057), .Z(n5778) );
  ANDN U5867 ( .A(n6058), .B(n6059), .Z(n6057) );
  XNOR U5868 ( .A(n6056), .B(n6060), .Z(n6058) );
  XOR U5869 ( .A(n5789), .B(n6061), .Z(n5782) );
  IV U5870 ( .A(n5788), .Z(n6061) );
  XNOR U5871 ( .A(n5785), .B(n6062), .Z(n5788) );
  XOR U5872 ( .A(n6063), .B(n6064), .Z(n5785) );
  ANDN U5873 ( .A(n6065), .B(n6066), .Z(n6064) );
  XNOR U5874 ( .A(n6063), .B(n6067), .Z(n6065) );
  XOR U5875 ( .A(n5796), .B(n6068), .Z(n5789) );
  IV U5876 ( .A(n5795), .Z(n6068) );
  XNOR U5877 ( .A(n5792), .B(n6069), .Z(n5795) );
  XOR U5878 ( .A(n6070), .B(n6071), .Z(n5792) );
  ANDN U5879 ( .A(n6072), .B(n6073), .Z(n6071) );
  XNOR U5880 ( .A(n6070), .B(n6074), .Z(n6072) );
  XOR U5881 ( .A(n5803), .B(n6075), .Z(n5796) );
  IV U5882 ( .A(n5802), .Z(n6075) );
  XNOR U5883 ( .A(n5799), .B(n6076), .Z(n5802) );
  XOR U5884 ( .A(n6077), .B(n6078), .Z(n5799) );
  ANDN U5885 ( .A(n6079), .B(n6080), .Z(n6078) );
  XNOR U5886 ( .A(n6077), .B(n6081), .Z(n6079) );
  XOR U5887 ( .A(n5810), .B(n6082), .Z(n5803) );
  IV U5888 ( .A(n5809), .Z(n6082) );
  XNOR U5889 ( .A(n5806), .B(n6083), .Z(n5809) );
  XOR U5890 ( .A(n6084), .B(n6085), .Z(n5806) );
  ANDN U5891 ( .A(n6086), .B(n6087), .Z(n6085) );
  XNOR U5892 ( .A(n6084), .B(n6088), .Z(n6086) );
  XOR U5893 ( .A(n5817), .B(n6089), .Z(n5810) );
  IV U5894 ( .A(n5816), .Z(n6089) );
  XNOR U5895 ( .A(n5813), .B(n6090), .Z(n5816) );
  XOR U5896 ( .A(n6091), .B(n6092), .Z(n5813) );
  ANDN U5897 ( .A(n6093), .B(n6094), .Z(n6092) );
  XNOR U5898 ( .A(n6091), .B(n6095), .Z(n6093) );
  XOR U5899 ( .A(n5824), .B(n6096), .Z(n5817) );
  IV U5900 ( .A(n5823), .Z(n6096) );
  XNOR U5901 ( .A(n5820), .B(n6097), .Z(n5823) );
  XOR U5902 ( .A(n6098), .B(n6099), .Z(n5820) );
  ANDN U5903 ( .A(n6100), .B(n6101), .Z(n6099) );
  XNOR U5904 ( .A(n6098), .B(n6102), .Z(n6100) );
  XOR U5905 ( .A(n5831), .B(n6103), .Z(n5824) );
  IV U5906 ( .A(n5830), .Z(n6103) );
  XNOR U5907 ( .A(n5827), .B(n6104), .Z(n5830) );
  XOR U5908 ( .A(n6105), .B(n6106), .Z(n5827) );
  ANDN U5909 ( .A(n6107), .B(n6108), .Z(n6106) );
  XNOR U5910 ( .A(n6105), .B(n6109), .Z(n6107) );
  XOR U5911 ( .A(n5838), .B(n6110), .Z(n5831) );
  IV U5912 ( .A(n5837), .Z(n6110) );
  XNOR U5913 ( .A(n5834), .B(n6111), .Z(n5837) );
  XOR U5914 ( .A(n6112), .B(n6113), .Z(n5834) );
  ANDN U5915 ( .A(n6114), .B(n6115), .Z(n6113) );
  XNOR U5916 ( .A(n6112), .B(n6116), .Z(n6114) );
  XOR U5917 ( .A(n5844), .B(n6117), .Z(n5838) );
  IV U5918 ( .A(n5843), .Z(n6117) );
  XNOR U5919 ( .A(n5840), .B(n6118), .Z(n5843) );
  XOR U5920 ( .A(n6119), .B(n6120), .Z(n5840) );
  ANDN U5921 ( .A(n6121), .B(n6122), .Z(n6120) );
  XNOR U5922 ( .A(n6119), .B(n6123), .Z(n6121) );
  XOR U5923 ( .A(n5850), .B(n6124), .Z(n5844) );
  IV U5924 ( .A(n5849), .Z(n6124) );
  XNOR U5925 ( .A(n5846), .B(n6111), .Z(n5849) );
  AND U5926 ( .A(n6688), .B(n5561), .Z(n6111) );
  XOR U5927 ( .A(n6125), .B(n6126), .Z(n5846) );
  ANDN U5928 ( .A(n6127), .B(n6128), .Z(n6126) );
  XNOR U5929 ( .A(n6125), .B(n6129), .Z(n6127) );
  XOR U5930 ( .A(n5856), .B(n6130), .Z(n5850) );
  IV U5931 ( .A(n5855), .Z(n6130) );
  XNOR U5932 ( .A(n5852), .B(n6104), .Z(n5855) );
  AND U5933 ( .A(n7241), .B(n5030), .Z(n6104) );
  XOR U5934 ( .A(n6131), .B(n6132), .Z(n5852) );
  ANDN U5935 ( .A(n6133), .B(n6134), .Z(n6132) );
  XNOR U5936 ( .A(n6131), .B(n6135), .Z(n6133) );
  XOR U5937 ( .A(n5862), .B(n6136), .Z(n5856) );
  IV U5938 ( .A(n5861), .Z(n6136) );
  XNOR U5939 ( .A(n5858), .B(n6097), .Z(n5861) );
  AND U5940 ( .A(n7770), .B(n4525), .Z(n6097) );
  XOR U5941 ( .A(n6137), .B(n6138), .Z(n5858) );
  ANDN U5942 ( .A(n6139), .B(n6140), .Z(n6138) );
  XNOR U5943 ( .A(n6137), .B(n6141), .Z(n6139) );
  XOR U5944 ( .A(n5868), .B(n6142), .Z(n5862) );
  IV U5945 ( .A(n5867), .Z(n6142) );
  XNOR U5946 ( .A(n5864), .B(n6090), .Z(n5867) );
  AND U5947 ( .A(n8272), .B(n4046), .Z(n6090) );
  XOR U5948 ( .A(n6143), .B(n6144), .Z(n5864) );
  ANDN U5949 ( .A(n6145), .B(n6146), .Z(n6144) );
  XNOR U5950 ( .A(n6143), .B(n6147), .Z(n6145) );
  XOR U5951 ( .A(n5874), .B(n6148), .Z(n5868) );
  IV U5952 ( .A(n5873), .Z(n6148) );
  XNOR U5953 ( .A(n5870), .B(n6083), .Z(n5873) );
  AND U5954 ( .A(n8748), .B(n3593), .Z(n6083) );
  XOR U5955 ( .A(n6149), .B(n6150), .Z(n5870) );
  ANDN U5956 ( .A(n6151), .B(n6152), .Z(n6150) );
  XNOR U5957 ( .A(n6149), .B(n6153), .Z(n6151) );
  XOR U5958 ( .A(n5880), .B(n6154), .Z(n5874) );
  IV U5959 ( .A(n5879), .Z(n6154) );
  XNOR U5960 ( .A(n5876), .B(n6076), .Z(n5879) );
  AND U5961 ( .A(n9198), .B(n3166), .Z(n6076) );
  XOR U5962 ( .A(n6155), .B(n6156), .Z(n5876) );
  ANDN U5963 ( .A(n6157), .B(n6158), .Z(n6156) );
  XNOR U5964 ( .A(n6155), .B(n6159), .Z(n6157) );
  XOR U5965 ( .A(n5886), .B(n6160), .Z(n5880) );
  IV U5966 ( .A(n5885), .Z(n6160) );
  XNOR U5967 ( .A(n5882), .B(n6069), .Z(n5885) );
  AND U5968 ( .A(n9621), .B(n2765), .Z(n6069) );
  XOR U5969 ( .A(n6161), .B(n6162), .Z(n5882) );
  ANDN U5970 ( .A(n6163), .B(n6164), .Z(n6162) );
  XNOR U5971 ( .A(n6161), .B(n6165), .Z(n6163) );
  XOR U5972 ( .A(n5892), .B(n6166), .Z(n5886) );
  IV U5973 ( .A(n5891), .Z(n6166) );
  XNOR U5974 ( .A(n5888), .B(n6062), .Z(n5891) );
  AND U5975 ( .A(n10017), .B(n2396), .Z(n6062) );
  XOR U5976 ( .A(n6167), .B(n6168), .Z(n5888) );
  ANDN U5977 ( .A(n6169), .B(n6170), .Z(n6168) );
  XNOR U5978 ( .A(n6167), .B(n6171), .Z(n6169) );
  XOR U5979 ( .A(n5898), .B(n6172), .Z(n5892) );
  IV U5980 ( .A(n5897), .Z(n6172) );
  XNOR U5981 ( .A(n5894), .B(n6055), .Z(n5897) );
  AND U5982 ( .A(n10387), .B(n2053), .Z(n6055) );
  XOR U5983 ( .A(n6173), .B(n6174), .Z(n5894) );
  ANDN U5984 ( .A(n6175), .B(n6176), .Z(n6174) );
  XNOR U5985 ( .A(n6173), .B(n6177), .Z(n6175) );
  XOR U5986 ( .A(n5904), .B(n6178), .Z(n5898) );
  IV U5987 ( .A(n5903), .Z(n6178) );
  XNOR U5988 ( .A(n5900), .B(n6048), .Z(n5903) );
  AND U5989 ( .A(n10731), .B(n1737), .Z(n6048) );
  XOR U5990 ( .A(n6179), .B(n6180), .Z(n5900) );
  ANDN U5991 ( .A(n6181), .B(n6182), .Z(n6180) );
  XNOR U5992 ( .A(n6179), .B(n6183), .Z(n6181) );
  XOR U5993 ( .A(n5910), .B(n6184), .Z(n5904) );
  IV U5994 ( .A(n5909), .Z(n6184) );
  XNOR U5995 ( .A(n5906), .B(n6041), .Z(n5909) );
  AND U5996 ( .A(n11049), .B(n1448), .Z(n6041) );
  XOR U5997 ( .A(n6185), .B(n6186), .Z(n5906) );
  ANDN U5998 ( .A(n6187), .B(n6188), .Z(n6186) );
  XNOR U5999 ( .A(n6185), .B(n6189), .Z(n6187) );
  XOR U6000 ( .A(n5916), .B(n6190), .Z(n5910) );
  IV U6001 ( .A(n5915), .Z(n6190) );
  XNOR U6002 ( .A(n5912), .B(n6034), .Z(n5915) );
  AND U6003 ( .A(n11341), .B(n1185), .Z(n6034) );
  XOR U6004 ( .A(n6191), .B(n6192), .Z(n5912) );
  ANDN U6005 ( .A(n6193), .B(n6194), .Z(n6192) );
  XNOR U6006 ( .A(n6191), .B(n6195), .Z(n6193) );
  XOR U6007 ( .A(n5922), .B(n6196), .Z(n5916) );
  IV U6008 ( .A(n5921), .Z(n6196) );
  XNOR U6009 ( .A(n5918), .B(n6027), .Z(n5921) );
  AND U6010 ( .A(n11607), .B(n948), .Z(n6027) );
  XOR U6011 ( .A(n6197), .B(n6198), .Z(n5918) );
  ANDN U6012 ( .A(n6199), .B(n6200), .Z(n6198) );
  XNOR U6013 ( .A(n6197), .B(n6201), .Z(n6199) );
  XOR U6014 ( .A(n5928), .B(n6202), .Z(n5922) );
  IV U6015 ( .A(n5927), .Z(n6202) );
  XNOR U6016 ( .A(n5924), .B(n6020), .Z(n5927) );
  AND U6017 ( .A(n11869), .B(n736), .Z(n6020) );
  XOR U6018 ( .A(n6203), .B(n6204), .Z(n5924) );
  ANDN U6019 ( .A(n6205), .B(n6206), .Z(n6204) );
  XNOR U6020 ( .A(n6203), .B(n6207), .Z(n6205) );
  XOR U6021 ( .A(n5934), .B(n6208), .Z(n5928) );
  IV U6022 ( .A(n5933), .Z(n6208) );
  XNOR U6023 ( .A(n5930), .B(n6013), .Z(n5933) );
  AND U6024 ( .A(n12128), .B(n552), .Z(n6013) );
  XOR U6025 ( .A(n6209), .B(n6210), .Z(n5930) );
  ANDN U6026 ( .A(n6211), .B(n6212), .Z(n6210) );
  XNOR U6027 ( .A(n6209), .B(n6213), .Z(n6211) );
  XOR U6028 ( .A(n5940), .B(n6214), .Z(n5934) );
  IV U6029 ( .A(n5939), .Z(n6214) );
  XNOR U6030 ( .A(n5936), .B(n6006), .Z(n5939) );
  AND U6031 ( .A(n12387), .B(n395), .Z(n6006) );
  XOR U6032 ( .A(n6215), .B(n6216), .Z(n5936) );
  ANDN U6033 ( .A(n6217), .B(n6218), .Z(n6216) );
  XNOR U6034 ( .A(n6215), .B(n6219), .Z(n6217) );
  XOR U6035 ( .A(n5946), .B(n6220), .Z(n5940) );
  IV U6036 ( .A(n5945), .Z(n6220) );
  XNOR U6037 ( .A(n5942), .B(n5999), .Z(n5945) );
  AND U6038 ( .A(n12644), .B(n264), .Z(n5999) );
  XOR U6039 ( .A(n6221), .B(n6222), .Z(n5942) );
  ANDN U6040 ( .A(n6223), .B(n6224), .Z(n6222) );
  XNOR U6041 ( .A(n6221), .B(n6225), .Z(n6223) );
  XOR U6042 ( .A(n5952), .B(n6226), .Z(n5946) );
  IV U6043 ( .A(n5951), .Z(n6226) );
  XNOR U6044 ( .A(n5948), .B(n5992), .Z(n5951) );
  AND U6045 ( .A(n12880), .B(n159), .Z(n5992) );
  XOR U6046 ( .A(n6227), .B(n6228), .Z(n5948) );
  ANDN U6047 ( .A(n6229), .B(n6230), .Z(n6228) );
  XNOR U6048 ( .A(n6227), .B(n6231), .Z(n6229) );
  XOR U6049 ( .A(n5959), .B(n6232), .Z(n5952) );
  IV U6050 ( .A(n5958), .Z(n6232) );
  XNOR U6051 ( .A(n5955), .B(n5985), .Z(n5958) );
  AND U6052 ( .A(n13070), .B(n80), .Z(n5985) );
  XOR U6053 ( .A(n6233), .B(n6234), .Z(n5955) );
  ANDN U6054 ( .A(n6235), .B(n6236), .Z(n6234) );
  XNOR U6055 ( .A(n6233), .B(n6237), .Z(n6235) );
  XOR U6056 ( .A(n5964), .B(n6238), .Z(n5959) );
  IV U6057 ( .A(n5963), .Z(n6238) );
  XNOR U6058 ( .A(n5960), .B(n6239), .Z(n5963) );
  AND U6059 ( .A(n42), .B(n13207), .Z(n6239) );
  XOR U6060 ( .A(n6240), .B(n6241), .Z(n5960) );
  ANDN U6061 ( .A(n6242), .B(n6243), .Z(n6241) );
  XOR U6062 ( .A(n6240), .B(n6244), .Z(n6242) );
  XNOR U6063 ( .A(n6245), .B(n6246), .Z(n5964) );
  ANDN U6064 ( .A(n6245), .B(n6247), .Z(n6246) );
  XNOR U6065 ( .A(n5973), .B(n5965), .Z(n5983) );
  XOR U6066 ( .A(n6248), .B(n6249), .Z(n5965) );
  AND U6067 ( .A(n6250), .B(n6251), .Z(n6249) );
  XNOR U6068 ( .A(n6252), .B(n6248), .Z(n6251) );
  XOR U6069 ( .A(n5971), .B(n6253), .Z(n5973) );
  ANDN U6070 ( .A(n13207), .B(n43), .Z(n6253) );
  XOR U6071 ( .A(n6254), .B(n6255), .Z(n5971) );
  NAND U6072 ( .A(n6256), .B(n6257), .Z(n6254) );
  XOR U6073 ( .A(n6255), .B(n6258), .Z(n6256) );
  XOR U6074 ( .A(n5969), .B(n5979), .Z(n5982) );
  XOR U6075 ( .A(n6259), .B(n6260), .Z(n5969) );
  IV U6076 ( .A(n6261), .Z(n6260) );
  XOR U6077 ( .A(n6262), .B(n6263), .Z(n5979) );
  AND U6078 ( .A(n6262), .B(n6264), .Z(n6263) );
  XOR U6079 ( .A(n6265), .B(n6250), .Z(n6264) );
  XOR U6080 ( .A(n6266), .B(n6258), .Z(n6250) );
  XOR U6081 ( .A(n5990), .B(n6267), .Z(n6258) );
  IV U6082 ( .A(n5989), .Z(n6267) );
  XNOR U6083 ( .A(n5986), .B(n6268), .Z(n5989) );
  XOR U6084 ( .A(n6269), .B(n6270), .Z(n5986) );
  NANDN U6085 ( .B(n6271), .A(n6272), .Z(n6269) );
  XOR U6086 ( .A(n6270), .B(n6273), .Z(n6272) );
  XOR U6087 ( .A(n5997), .B(n6274), .Z(n5990) );
  IV U6088 ( .A(n5996), .Z(n6274) );
  XNOR U6089 ( .A(n5993), .B(n6275), .Z(n5996) );
  XOR U6090 ( .A(n6276), .B(n6277), .Z(n5993) );
  ANDN U6091 ( .A(n6278), .B(n6279), .Z(n6277) );
  XNOR U6092 ( .A(n6276), .B(n6280), .Z(n6278) );
  XOR U6093 ( .A(n6004), .B(n6281), .Z(n5997) );
  IV U6094 ( .A(n6003), .Z(n6281) );
  XNOR U6095 ( .A(n6000), .B(n6282), .Z(n6003) );
  XOR U6096 ( .A(n6283), .B(n6284), .Z(n6000) );
  ANDN U6097 ( .A(n6285), .B(n6286), .Z(n6284) );
  XNOR U6098 ( .A(n6283), .B(n6287), .Z(n6285) );
  XOR U6099 ( .A(n6011), .B(n6288), .Z(n6004) );
  IV U6100 ( .A(n6010), .Z(n6288) );
  XNOR U6101 ( .A(n6007), .B(n6289), .Z(n6010) );
  XOR U6102 ( .A(n6290), .B(n6291), .Z(n6007) );
  ANDN U6103 ( .A(n6292), .B(n6293), .Z(n6291) );
  XNOR U6104 ( .A(n6290), .B(n6294), .Z(n6292) );
  XOR U6105 ( .A(n6018), .B(n6295), .Z(n6011) );
  IV U6106 ( .A(n6017), .Z(n6295) );
  XNOR U6107 ( .A(n6014), .B(n6296), .Z(n6017) );
  XOR U6108 ( .A(n6297), .B(n6298), .Z(n6014) );
  ANDN U6109 ( .A(n6299), .B(n6300), .Z(n6298) );
  XNOR U6110 ( .A(n6297), .B(n6301), .Z(n6299) );
  XOR U6111 ( .A(n6025), .B(n6302), .Z(n6018) );
  IV U6112 ( .A(n6024), .Z(n6302) );
  XNOR U6113 ( .A(n6021), .B(n6303), .Z(n6024) );
  XOR U6114 ( .A(n6304), .B(n6305), .Z(n6021) );
  ANDN U6115 ( .A(n6306), .B(n6307), .Z(n6305) );
  XNOR U6116 ( .A(n6304), .B(n6308), .Z(n6306) );
  XOR U6117 ( .A(n6032), .B(n6309), .Z(n6025) );
  IV U6118 ( .A(n6031), .Z(n6309) );
  XNOR U6119 ( .A(n6028), .B(n6310), .Z(n6031) );
  XOR U6120 ( .A(n6311), .B(n6312), .Z(n6028) );
  ANDN U6121 ( .A(n6313), .B(n6314), .Z(n6312) );
  XNOR U6122 ( .A(n6311), .B(n6315), .Z(n6313) );
  XOR U6123 ( .A(n6039), .B(n6316), .Z(n6032) );
  IV U6124 ( .A(n6038), .Z(n6316) );
  XNOR U6125 ( .A(n6035), .B(n6317), .Z(n6038) );
  XOR U6126 ( .A(n6318), .B(n6319), .Z(n6035) );
  ANDN U6127 ( .A(n6320), .B(n6321), .Z(n6319) );
  XNOR U6128 ( .A(n6318), .B(n6322), .Z(n6320) );
  XOR U6129 ( .A(n6046), .B(n6323), .Z(n6039) );
  IV U6130 ( .A(n6045), .Z(n6323) );
  XNOR U6131 ( .A(n6042), .B(n6324), .Z(n6045) );
  XOR U6132 ( .A(n6325), .B(n6326), .Z(n6042) );
  ANDN U6133 ( .A(n6327), .B(n6328), .Z(n6326) );
  XNOR U6134 ( .A(n6325), .B(n6329), .Z(n6327) );
  XOR U6135 ( .A(n6053), .B(n6330), .Z(n6046) );
  IV U6136 ( .A(n6052), .Z(n6330) );
  XNOR U6137 ( .A(n6049), .B(n6331), .Z(n6052) );
  XOR U6138 ( .A(n6332), .B(n6333), .Z(n6049) );
  ANDN U6139 ( .A(n6334), .B(n6335), .Z(n6333) );
  XNOR U6140 ( .A(n6332), .B(n6336), .Z(n6334) );
  XOR U6141 ( .A(n6060), .B(n6337), .Z(n6053) );
  IV U6142 ( .A(n6059), .Z(n6337) );
  XNOR U6143 ( .A(n6056), .B(n6338), .Z(n6059) );
  XOR U6144 ( .A(n6339), .B(n6340), .Z(n6056) );
  ANDN U6145 ( .A(n6341), .B(n6342), .Z(n6340) );
  XNOR U6146 ( .A(n6339), .B(n6343), .Z(n6341) );
  XOR U6147 ( .A(n6067), .B(n6344), .Z(n6060) );
  IV U6148 ( .A(n6066), .Z(n6344) );
  XNOR U6149 ( .A(n6063), .B(n6345), .Z(n6066) );
  XOR U6150 ( .A(n6346), .B(n6347), .Z(n6063) );
  ANDN U6151 ( .A(n6348), .B(n6349), .Z(n6347) );
  XNOR U6152 ( .A(n6346), .B(n6350), .Z(n6348) );
  XOR U6153 ( .A(n6074), .B(n6351), .Z(n6067) );
  IV U6154 ( .A(n6073), .Z(n6351) );
  XNOR U6155 ( .A(n6070), .B(n6352), .Z(n6073) );
  XOR U6156 ( .A(n6353), .B(n6354), .Z(n6070) );
  ANDN U6157 ( .A(n6355), .B(n6356), .Z(n6354) );
  XNOR U6158 ( .A(n6353), .B(n6357), .Z(n6355) );
  XOR U6159 ( .A(n6081), .B(n6358), .Z(n6074) );
  IV U6160 ( .A(n6080), .Z(n6358) );
  XNOR U6161 ( .A(n6077), .B(n6359), .Z(n6080) );
  XOR U6162 ( .A(n6360), .B(n6361), .Z(n6077) );
  ANDN U6163 ( .A(n6362), .B(n6363), .Z(n6361) );
  XNOR U6164 ( .A(n6360), .B(n6364), .Z(n6362) );
  XOR U6165 ( .A(n6088), .B(n6365), .Z(n6081) );
  IV U6166 ( .A(n6087), .Z(n6365) );
  XNOR U6167 ( .A(n6084), .B(n6366), .Z(n6087) );
  XOR U6168 ( .A(n6367), .B(n6368), .Z(n6084) );
  ANDN U6169 ( .A(n6369), .B(n6370), .Z(n6368) );
  XNOR U6170 ( .A(n6367), .B(n6371), .Z(n6369) );
  XOR U6171 ( .A(n6095), .B(n6372), .Z(n6088) );
  IV U6172 ( .A(n6094), .Z(n6372) );
  XNOR U6173 ( .A(n6091), .B(n6373), .Z(n6094) );
  XOR U6174 ( .A(n6374), .B(n6375), .Z(n6091) );
  ANDN U6175 ( .A(n6376), .B(n6377), .Z(n6375) );
  XNOR U6176 ( .A(n6374), .B(n6378), .Z(n6376) );
  XOR U6177 ( .A(n6102), .B(n6379), .Z(n6095) );
  IV U6178 ( .A(n6101), .Z(n6379) );
  XNOR U6179 ( .A(n6098), .B(n6380), .Z(n6101) );
  XOR U6180 ( .A(n6381), .B(n6382), .Z(n6098) );
  ANDN U6181 ( .A(n6383), .B(n6384), .Z(n6382) );
  XNOR U6182 ( .A(n6381), .B(n6385), .Z(n6383) );
  XOR U6183 ( .A(n6109), .B(n6386), .Z(n6102) );
  IV U6184 ( .A(n6108), .Z(n6386) );
  XNOR U6185 ( .A(n6105), .B(n6387), .Z(n6108) );
  XOR U6186 ( .A(n6388), .B(n6389), .Z(n6105) );
  ANDN U6187 ( .A(n6390), .B(n6391), .Z(n6389) );
  XNOR U6188 ( .A(n6388), .B(n6392), .Z(n6390) );
  XOR U6189 ( .A(n6116), .B(n6393), .Z(n6109) );
  IV U6190 ( .A(n6115), .Z(n6393) );
  XNOR U6191 ( .A(n6112), .B(n6394), .Z(n6115) );
  XOR U6192 ( .A(n6395), .B(n6396), .Z(n6112) );
  ANDN U6193 ( .A(n6397), .B(n6398), .Z(n6396) );
  XNOR U6194 ( .A(n6395), .B(n6399), .Z(n6397) );
  XOR U6195 ( .A(n6123), .B(n6400), .Z(n6116) );
  IV U6196 ( .A(n6122), .Z(n6400) );
  XNOR U6197 ( .A(n6119), .B(n6401), .Z(n6122) );
  XOR U6198 ( .A(n6402), .B(n6403), .Z(n6119) );
  ANDN U6199 ( .A(n6404), .B(n6405), .Z(n6403) );
  XNOR U6200 ( .A(n6402), .B(n6406), .Z(n6404) );
  XOR U6201 ( .A(n6129), .B(n6407), .Z(n6123) );
  IV U6202 ( .A(n6128), .Z(n6407) );
  XNOR U6203 ( .A(n6125), .B(n6401), .Z(n6128) );
  AND U6204 ( .A(n6688), .B(n6118), .Z(n6401) );
  XOR U6205 ( .A(n6408), .B(n6409), .Z(n6125) );
  ANDN U6206 ( .A(n6410), .B(n6411), .Z(n6409) );
  XNOR U6207 ( .A(n6408), .B(n6412), .Z(n6410) );
  XOR U6208 ( .A(n6135), .B(n6413), .Z(n6129) );
  IV U6209 ( .A(n6134), .Z(n6413) );
  XNOR U6210 ( .A(n6131), .B(n6394), .Z(n6134) );
  AND U6211 ( .A(n7241), .B(n5561), .Z(n6394) );
  XOR U6212 ( .A(n6414), .B(n6415), .Z(n6131) );
  ANDN U6213 ( .A(n6416), .B(n6417), .Z(n6415) );
  XNOR U6214 ( .A(n6414), .B(n6418), .Z(n6416) );
  XOR U6215 ( .A(n6141), .B(n6419), .Z(n6135) );
  IV U6216 ( .A(n6140), .Z(n6419) );
  XNOR U6217 ( .A(n6137), .B(n6387), .Z(n6140) );
  AND U6218 ( .A(n7770), .B(n5030), .Z(n6387) );
  XOR U6219 ( .A(n6420), .B(n6421), .Z(n6137) );
  ANDN U6220 ( .A(n6422), .B(n6423), .Z(n6421) );
  XNOR U6221 ( .A(n6420), .B(n6424), .Z(n6422) );
  XOR U6222 ( .A(n6147), .B(n6425), .Z(n6141) );
  IV U6223 ( .A(n6146), .Z(n6425) );
  XNOR U6224 ( .A(n6143), .B(n6380), .Z(n6146) );
  AND U6225 ( .A(n8272), .B(n4525), .Z(n6380) );
  XOR U6226 ( .A(n6426), .B(n6427), .Z(n6143) );
  ANDN U6227 ( .A(n6428), .B(n6429), .Z(n6427) );
  XNOR U6228 ( .A(n6426), .B(n6430), .Z(n6428) );
  XOR U6229 ( .A(n6153), .B(n6431), .Z(n6147) );
  IV U6230 ( .A(n6152), .Z(n6431) );
  XNOR U6231 ( .A(n6149), .B(n6373), .Z(n6152) );
  AND U6232 ( .A(n8748), .B(n4046), .Z(n6373) );
  XOR U6233 ( .A(n6432), .B(n6433), .Z(n6149) );
  ANDN U6234 ( .A(n6434), .B(n6435), .Z(n6433) );
  XNOR U6235 ( .A(n6432), .B(n6436), .Z(n6434) );
  XOR U6236 ( .A(n6159), .B(n6437), .Z(n6153) );
  IV U6237 ( .A(n6158), .Z(n6437) );
  XNOR U6238 ( .A(n6155), .B(n6366), .Z(n6158) );
  AND U6239 ( .A(n9198), .B(n3593), .Z(n6366) );
  XOR U6240 ( .A(n6438), .B(n6439), .Z(n6155) );
  ANDN U6241 ( .A(n6440), .B(n6441), .Z(n6439) );
  XNOR U6242 ( .A(n6438), .B(n6442), .Z(n6440) );
  XOR U6243 ( .A(n6165), .B(n6443), .Z(n6159) );
  IV U6244 ( .A(n6164), .Z(n6443) );
  XNOR U6245 ( .A(n6161), .B(n6359), .Z(n6164) );
  AND U6246 ( .A(n9621), .B(n3166), .Z(n6359) );
  XOR U6247 ( .A(n6444), .B(n6445), .Z(n6161) );
  ANDN U6248 ( .A(n6446), .B(n6447), .Z(n6445) );
  XNOR U6249 ( .A(n6444), .B(n6448), .Z(n6446) );
  XOR U6250 ( .A(n6171), .B(n6449), .Z(n6165) );
  IV U6251 ( .A(n6170), .Z(n6449) );
  XNOR U6252 ( .A(n6167), .B(n6352), .Z(n6170) );
  AND U6253 ( .A(n10017), .B(n2765), .Z(n6352) );
  XOR U6254 ( .A(n6450), .B(n6451), .Z(n6167) );
  ANDN U6255 ( .A(n6452), .B(n6453), .Z(n6451) );
  XNOR U6256 ( .A(n6450), .B(n6454), .Z(n6452) );
  XOR U6257 ( .A(n6177), .B(n6455), .Z(n6171) );
  IV U6258 ( .A(n6176), .Z(n6455) );
  XNOR U6259 ( .A(n6173), .B(n6345), .Z(n6176) );
  AND U6260 ( .A(n10387), .B(n2396), .Z(n6345) );
  XOR U6261 ( .A(n6456), .B(n6457), .Z(n6173) );
  ANDN U6262 ( .A(n6458), .B(n6459), .Z(n6457) );
  XNOR U6263 ( .A(n6456), .B(n6460), .Z(n6458) );
  XOR U6264 ( .A(n6183), .B(n6461), .Z(n6177) );
  IV U6265 ( .A(n6182), .Z(n6461) );
  XNOR U6266 ( .A(n6179), .B(n6338), .Z(n6182) );
  AND U6267 ( .A(n10731), .B(n2053), .Z(n6338) );
  XOR U6268 ( .A(n6462), .B(n6463), .Z(n6179) );
  ANDN U6269 ( .A(n6464), .B(n6465), .Z(n6463) );
  XNOR U6270 ( .A(n6462), .B(n6466), .Z(n6464) );
  XOR U6271 ( .A(n6189), .B(n6467), .Z(n6183) );
  IV U6272 ( .A(n6188), .Z(n6467) );
  XNOR U6273 ( .A(n6185), .B(n6331), .Z(n6188) );
  AND U6274 ( .A(n11049), .B(n1737), .Z(n6331) );
  XOR U6275 ( .A(n6468), .B(n6469), .Z(n6185) );
  ANDN U6276 ( .A(n6470), .B(n6471), .Z(n6469) );
  XNOR U6277 ( .A(n6468), .B(n6472), .Z(n6470) );
  XOR U6278 ( .A(n6195), .B(n6473), .Z(n6189) );
  IV U6279 ( .A(n6194), .Z(n6473) );
  XNOR U6280 ( .A(n6191), .B(n6324), .Z(n6194) );
  AND U6281 ( .A(n11341), .B(n1448), .Z(n6324) );
  XOR U6282 ( .A(n6474), .B(n6475), .Z(n6191) );
  ANDN U6283 ( .A(n6476), .B(n6477), .Z(n6475) );
  XNOR U6284 ( .A(n6474), .B(n6478), .Z(n6476) );
  XOR U6285 ( .A(n6201), .B(n6479), .Z(n6195) );
  IV U6286 ( .A(n6200), .Z(n6479) );
  XNOR U6287 ( .A(n6197), .B(n6317), .Z(n6200) );
  AND U6288 ( .A(n11607), .B(n1185), .Z(n6317) );
  XOR U6289 ( .A(n6480), .B(n6481), .Z(n6197) );
  ANDN U6290 ( .A(n6482), .B(n6483), .Z(n6481) );
  XNOR U6291 ( .A(n6480), .B(n6484), .Z(n6482) );
  XOR U6292 ( .A(n6207), .B(n6485), .Z(n6201) );
  IV U6293 ( .A(n6206), .Z(n6485) );
  XNOR U6294 ( .A(n6203), .B(n6310), .Z(n6206) );
  AND U6295 ( .A(n11869), .B(n948), .Z(n6310) );
  XOR U6296 ( .A(n6486), .B(n6487), .Z(n6203) );
  ANDN U6297 ( .A(n6488), .B(n6489), .Z(n6487) );
  XNOR U6298 ( .A(n6486), .B(n6490), .Z(n6488) );
  XOR U6299 ( .A(n6213), .B(n6491), .Z(n6207) );
  IV U6300 ( .A(n6212), .Z(n6491) );
  XNOR U6301 ( .A(n6209), .B(n6303), .Z(n6212) );
  AND U6302 ( .A(n12128), .B(n736), .Z(n6303) );
  XOR U6303 ( .A(n6492), .B(n6493), .Z(n6209) );
  ANDN U6304 ( .A(n6494), .B(n6495), .Z(n6493) );
  XNOR U6305 ( .A(n6492), .B(n6496), .Z(n6494) );
  XOR U6306 ( .A(n6219), .B(n6497), .Z(n6213) );
  IV U6307 ( .A(n6218), .Z(n6497) );
  XNOR U6308 ( .A(n6215), .B(n6296), .Z(n6218) );
  AND U6309 ( .A(n12387), .B(n552), .Z(n6296) );
  XOR U6310 ( .A(n6498), .B(n6499), .Z(n6215) );
  ANDN U6311 ( .A(n6500), .B(n6501), .Z(n6499) );
  XNOR U6312 ( .A(n6498), .B(n6502), .Z(n6500) );
  XOR U6313 ( .A(n6225), .B(n6503), .Z(n6219) );
  IV U6314 ( .A(n6224), .Z(n6503) );
  XNOR U6315 ( .A(n6221), .B(n6289), .Z(n6224) );
  AND U6316 ( .A(n12644), .B(n395), .Z(n6289) );
  XOR U6317 ( .A(n6504), .B(n6505), .Z(n6221) );
  ANDN U6318 ( .A(n6506), .B(n6507), .Z(n6505) );
  XNOR U6319 ( .A(n6504), .B(n6508), .Z(n6506) );
  XOR U6320 ( .A(n6231), .B(n6509), .Z(n6225) );
  IV U6321 ( .A(n6230), .Z(n6509) );
  XNOR U6322 ( .A(n6227), .B(n6282), .Z(n6230) );
  AND U6323 ( .A(n12880), .B(n264), .Z(n6282) );
  XOR U6324 ( .A(n6510), .B(n6511), .Z(n6227) );
  ANDN U6325 ( .A(n6512), .B(n6513), .Z(n6511) );
  XNOR U6326 ( .A(n6510), .B(n6514), .Z(n6512) );
  XOR U6327 ( .A(n6237), .B(n6515), .Z(n6231) );
  IV U6328 ( .A(n6236), .Z(n6515) );
  XNOR U6329 ( .A(n6233), .B(n6275), .Z(n6236) );
  AND U6330 ( .A(n13070), .B(n159), .Z(n6275) );
  XOR U6331 ( .A(n6516), .B(n6517), .Z(n6233) );
  ANDN U6332 ( .A(n6518), .B(n6519), .Z(n6517) );
  XNOR U6333 ( .A(n6516), .B(n6520), .Z(n6518) );
  XOR U6334 ( .A(n6244), .B(n6243), .Z(n6237) );
  XNOR U6335 ( .A(n6240), .B(n6268), .Z(n6243) );
  AND U6336 ( .A(n13207), .B(n80), .Z(n6268) );
  XOR U6337 ( .A(n6521), .B(n6522), .Z(n6240) );
  ANDN U6338 ( .A(n6523), .B(n6524), .Z(n6522) );
  XNOR U6339 ( .A(n6521), .B(n6525), .Z(n6523) );
  IV U6340 ( .A(n6247), .Z(n6244) );
  XNOR U6341 ( .A(n6245), .B(n6526), .Z(n6247) );
  AND U6342 ( .A(n42), .B(n6527), .Z(n6526) );
  XOR U6343 ( .A(n6528), .B(n6529), .Z(n6245) );
  ANDN U6344 ( .A(n6530), .B(n6531), .Z(n6529) );
  XNOR U6345 ( .A(n6532), .B(n6528), .Z(n6530) );
  XNOR U6346 ( .A(n6257), .B(n6248), .Z(n6266) );
  XNOR U6347 ( .A(n6533), .B(n6534), .Z(n6248) );
  AND U6348 ( .A(n6535), .B(n6536), .Z(n6534) );
  XOR U6349 ( .A(n6537), .B(n6533), .Z(n6536) );
  XOR U6350 ( .A(n6538), .B(n6255), .Z(n6257) );
  OR U6351 ( .A(n6539), .B(n6540), .Z(n6255) );
  OR U6352 ( .A(n43), .B(n6541), .Z(n6538) );
  XOR U6353 ( .A(n6252), .B(n6262), .Z(n6265) );
  XOR U6354 ( .A(n6542), .B(n6543), .Z(n6252) );
  IV U6355 ( .A(n6544), .Z(n6543) );
  XOR U6356 ( .A(n6545), .B(n6546), .Z(n6262) );
  AND U6357 ( .A(n6545), .B(n6547), .Z(n6546) );
  XOR U6358 ( .A(n6548), .B(n6535), .Z(n6547) );
  XOR U6359 ( .A(n6549), .B(n6540), .Z(n6535) );
  XOR U6360 ( .A(n6273), .B(n6550), .Z(n6540) );
  IV U6361 ( .A(n6271), .Z(n6550) );
  XNOR U6362 ( .A(n6551), .B(n6270), .Z(n6271) );
  OR U6363 ( .A(n6552), .B(n6553), .Z(n6270) );
  NANDN U6364 ( .B(n6541), .A(n80), .Z(n6551) );
  XOR U6365 ( .A(n6280), .B(n6554), .Z(n6273) );
  IV U6366 ( .A(n6279), .Z(n6554) );
  XNOR U6367 ( .A(n6276), .B(n6555), .Z(n6279) );
  XOR U6368 ( .A(n6556), .B(n6557), .Z(n6276) );
  NANDN U6369 ( .B(n6558), .A(n6559), .Z(n6556) );
  XOR U6370 ( .A(n6557), .B(n6560), .Z(n6559) );
  XOR U6371 ( .A(n6287), .B(n6561), .Z(n6280) );
  IV U6372 ( .A(n6286), .Z(n6561) );
  XNOR U6373 ( .A(n6283), .B(n6562), .Z(n6286) );
  XOR U6374 ( .A(n6563), .B(n6564), .Z(n6283) );
  ANDN U6375 ( .A(n6565), .B(n6566), .Z(n6564) );
  XNOR U6376 ( .A(n6563), .B(n6567), .Z(n6565) );
  XOR U6377 ( .A(n6294), .B(n6568), .Z(n6287) );
  IV U6378 ( .A(n6293), .Z(n6568) );
  XNOR U6379 ( .A(n6290), .B(n6569), .Z(n6293) );
  XOR U6380 ( .A(n6570), .B(n6571), .Z(n6290) );
  ANDN U6381 ( .A(n6572), .B(n6573), .Z(n6571) );
  XNOR U6382 ( .A(n6570), .B(n6574), .Z(n6572) );
  XOR U6383 ( .A(n6301), .B(n6575), .Z(n6294) );
  IV U6384 ( .A(n6300), .Z(n6575) );
  XNOR U6385 ( .A(n6297), .B(n6576), .Z(n6300) );
  XOR U6386 ( .A(n6577), .B(n6578), .Z(n6297) );
  ANDN U6387 ( .A(n6579), .B(n6580), .Z(n6578) );
  XNOR U6388 ( .A(n6577), .B(n6581), .Z(n6579) );
  XOR U6389 ( .A(n6308), .B(n6582), .Z(n6301) );
  IV U6390 ( .A(n6307), .Z(n6582) );
  XNOR U6391 ( .A(n6304), .B(n6583), .Z(n6307) );
  XOR U6392 ( .A(n6584), .B(n6585), .Z(n6304) );
  ANDN U6393 ( .A(n6586), .B(n6587), .Z(n6585) );
  XNOR U6394 ( .A(n6584), .B(n6588), .Z(n6586) );
  XOR U6395 ( .A(n6315), .B(n6589), .Z(n6308) );
  IV U6396 ( .A(n6314), .Z(n6589) );
  XNOR U6397 ( .A(n6311), .B(n6590), .Z(n6314) );
  XOR U6398 ( .A(n6591), .B(n6592), .Z(n6311) );
  ANDN U6399 ( .A(n6593), .B(n6594), .Z(n6592) );
  XNOR U6400 ( .A(n6591), .B(n6595), .Z(n6593) );
  XOR U6401 ( .A(n6322), .B(n6596), .Z(n6315) );
  IV U6402 ( .A(n6321), .Z(n6596) );
  XNOR U6403 ( .A(n6318), .B(n6597), .Z(n6321) );
  XOR U6404 ( .A(n6598), .B(n6599), .Z(n6318) );
  ANDN U6405 ( .A(n6600), .B(n6601), .Z(n6599) );
  XNOR U6406 ( .A(n6598), .B(n6602), .Z(n6600) );
  XOR U6407 ( .A(n6329), .B(n6603), .Z(n6322) );
  IV U6408 ( .A(n6328), .Z(n6603) );
  XNOR U6409 ( .A(n6325), .B(n6604), .Z(n6328) );
  XOR U6410 ( .A(n6605), .B(n6606), .Z(n6325) );
  ANDN U6411 ( .A(n6607), .B(n6608), .Z(n6606) );
  XNOR U6412 ( .A(n6605), .B(n6609), .Z(n6607) );
  XOR U6413 ( .A(n6336), .B(n6610), .Z(n6329) );
  IV U6414 ( .A(n6335), .Z(n6610) );
  XNOR U6415 ( .A(n6332), .B(n6611), .Z(n6335) );
  XOR U6416 ( .A(n6612), .B(n6613), .Z(n6332) );
  ANDN U6417 ( .A(n6614), .B(n6615), .Z(n6613) );
  XNOR U6418 ( .A(n6612), .B(n6616), .Z(n6614) );
  XOR U6419 ( .A(n6343), .B(n6617), .Z(n6336) );
  IV U6420 ( .A(n6342), .Z(n6617) );
  XNOR U6421 ( .A(n6339), .B(n6618), .Z(n6342) );
  XOR U6422 ( .A(n6619), .B(n6620), .Z(n6339) );
  ANDN U6423 ( .A(n6621), .B(n6622), .Z(n6620) );
  XNOR U6424 ( .A(n6619), .B(n6623), .Z(n6621) );
  XOR U6425 ( .A(n6350), .B(n6624), .Z(n6343) );
  IV U6426 ( .A(n6349), .Z(n6624) );
  XNOR U6427 ( .A(n6346), .B(n6625), .Z(n6349) );
  XOR U6428 ( .A(n6626), .B(n6627), .Z(n6346) );
  ANDN U6429 ( .A(n6628), .B(n6629), .Z(n6627) );
  XNOR U6430 ( .A(n6626), .B(n6630), .Z(n6628) );
  XOR U6431 ( .A(n6357), .B(n6631), .Z(n6350) );
  IV U6432 ( .A(n6356), .Z(n6631) );
  XNOR U6433 ( .A(n6353), .B(n6632), .Z(n6356) );
  XOR U6434 ( .A(n6633), .B(n6634), .Z(n6353) );
  ANDN U6435 ( .A(n6635), .B(n6636), .Z(n6634) );
  XNOR U6436 ( .A(n6633), .B(n6637), .Z(n6635) );
  XOR U6437 ( .A(n6364), .B(n6638), .Z(n6357) );
  IV U6438 ( .A(n6363), .Z(n6638) );
  XNOR U6439 ( .A(n6360), .B(n6639), .Z(n6363) );
  XOR U6440 ( .A(n6640), .B(n6641), .Z(n6360) );
  ANDN U6441 ( .A(n6642), .B(n6643), .Z(n6641) );
  XNOR U6442 ( .A(n6640), .B(n6644), .Z(n6642) );
  XOR U6443 ( .A(n6371), .B(n6645), .Z(n6364) );
  IV U6444 ( .A(n6370), .Z(n6645) );
  XNOR U6445 ( .A(n6367), .B(n6646), .Z(n6370) );
  XOR U6446 ( .A(n6647), .B(n6648), .Z(n6367) );
  ANDN U6447 ( .A(n6649), .B(n6650), .Z(n6648) );
  XNOR U6448 ( .A(n6647), .B(n6651), .Z(n6649) );
  XOR U6449 ( .A(n6378), .B(n6652), .Z(n6371) );
  IV U6450 ( .A(n6377), .Z(n6652) );
  XNOR U6451 ( .A(n6374), .B(n6653), .Z(n6377) );
  XOR U6452 ( .A(n6654), .B(n6655), .Z(n6374) );
  ANDN U6453 ( .A(n6656), .B(n6657), .Z(n6655) );
  XNOR U6454 ( .A(n6654), .B(n6658), .Z(n6656) );
  XOR U6455 ( .A(n6385), .B(n6659), .Z(n6378) );
  IV U6456 ( .A(n6384), .Z(n6659) );
  XNOR U6457 ( .A(n6381), .B(n6660), .Z(n6384) );
  XOR U6458 ( .A(n6661), .B(n6662), .Z(n6381) );
  ANDN U6459 ( .A(n6663), .B(n6664), .Z(n6662) );
  XNOR U6460 ( .A(n6661), .B(n6665), .Z(n6663) );
  XOR U6461 ( .A(n6392), .B(n6666), .Z(n6385) );
  IV U6462 ( .A(n6391), .Z(n6666) );
  XNOR U6463 ( .A(n6388), .B(n6667), .Z(n6391) );
  XOR U6464 ( .A(n6668), .B(n6669), .Z(n6388) );
  ANDN U6465 ( .A(n6670), .B(n6671), .Z(n6669) );
  XNOR U6466 ( .A(n6668), .B(n6672), .Z(n6670) );
  XOR U6467 ( .A(n6399), .B(n6673), .Z(n6392) );
  IV U6468 ( .A(n6398), .Z(n6673) );
  XNOR U6469 ( .A(n6395), .B(n6674), .Z(n6398) );
  XOR U6470 ( .A(n6675), .B(n6676), .Z(n6395) );
  ANDN U6471 ( .A(n6677), .B(n6678), .Z(n6676) );
  XNOR U6472 ( .A(n6675), .B(n6679), .Z(n6677) );
  XOR U6473 ( .A(n6406), .B(n6680), .Z(n6399) );
  IV U6474 ( .A(n6405), .Z(n6680) );
  XNOR U6475 ( .A(n6402), .B(n6681), .Z(n6405) );
  XOR U6476 ( .A(n6682), .B(n6683), .Z(n6402) );
  ANDN U6477 ( .A(n6684), .B(n6685), .Z(n6683) );
  XNOR U6478 ( .A(n6682), .B(n6686), .Z(n6684) );
  XOR U6479 ( .A(n6412), .B(n6687), .Z(n6406) );
  IV U6480 ( .A(n6411), .Z(n6687) );
  XNOR U6481 ( .A(n6408), .B(n6688), .Z(n6411) );
  XOR U6482 ( .A(n6689), .B(n6690), .Z(n6408) );
  ANDN U6483 ( .A(n6691), .B(n6692), .Z(n6690) );
  XNOR U6484 ( .A(n6689), .B(n6693), .Z(n6691) );
  XOR U6485 ( .A(n6418), .B(n6694), .Z(n6412) );
  IV U6486 ( .A(n6417), .Z(n6694) );
  XNOR U6487 ( .A(n6414), .B(n6681), .Z(n6417) );
  AND U6488 ( .A(n7241), .B(n6118), .Z(n6681) );
  XOR U6489 ( .A(n6695), .B(n6696), .Z(n6414) );
  ANDN U6490 ( .A(n6697), .B(n6698), .Z(n6696) );
  XNOR U6491 ( .A(n6695), .B(n6699), .Z(n6697) );
  XOR U6492 ( .A(n6424), .B(n6700), .Z(n6418) );
  IV U6493 ( .A(n6423), .Z(n6700) );
  XNOR U6494 ( .A(n6420), .B(n6674), .Z(n6423) );
  AND U6495 ( .A(n7770), .B(n5561), .Z(n6674) );
  XOR U6496 ( .A(n6701), .B(n6702), .Z(n6420) );
  ANDN U6497 ( .A(n6703), .B(n6704), .Z(n6702) );
  XNOR U6498 ( .A(n6701), .B(n6705), .Z(n6703) );
  XOR U6499 ( .A(n6430), .B(n6706), .Z(n6424) );
  IV U6500 ( .A(n6429), .Z(n6706) );
  XNOR U6501 ( .A(n6426), .B(n6667), .Z(n6429) );
  AND U6502 ( .A(n8272), .B(n5030), .Z(n6667) );
  XOR U6503 ( .A(n6707), .B(n6708), .Z(n6426) );
  ANDN U6504 ( .A(n6709), .B(n6710), .Z(n6708) );
  XNOR U6505 ( .A(n6707), .B(n6711), .Z(n6709) );
  XOR U6506 ( .A(n6436), .B(n6712), .Z(n6430) );
  IV U6507 ( .A(n6435), .Z(n6712) );
  XNOR U6508 ( .A(n6432), .B(n6660), .Z(n6435) );
  AND U6509 ( .A(n8748), .B(n4525), .Z(n6660) );
  XOR U6510 ( .A(n6713), .B(n6714), .Z(n6432) );
  ANDN U6511 ( .A(n6715), .B(n6716), .Z(n6714) );
  XNOR U6512 ( .A(n6713), .B(n6717), .Z(n6715) );
  XOR U6513 ( .A(n6442), .B(n6718), .Z(n6436) );
  IV U6514 ( .A(n6441), .Z(n6718) );
  XNOR U6515 ( .A(n6438), .B(n6653), .Z(n6441) );
  AND U6516 ( .A(n9198), .B(n4046), .Z(n6653) );
  XOR U6517 ( .A(n6719), .B(n6720), .Z(n6438) );
  ANDN U6518 ( .A(n6721), .B(n6722), .Z(n6720) );
  XNOR U6519 ( .A(n6719), .B(n6723), .Z(n6721) );
  XOR U6520 ( .A(n6448), .B(n6724), .Z(n6442) );
  IV U6521 ( .A(n6447), .Z(n6724) );
  XNOR U6522 ( .A(n6444), .B(n6646), .Z(n6447) );
  AND U6523 ( .A(n9621), .B(n3593), .Z(n6646) );
  XOR U6524 ( .A(n6725), .B(n6726), .Z(n6444) );
  ANDN U6525 ( .A(n6727), .B(n6728), .Z(n6726) );
  XNOR U6526 ( .A(n6725), .B(n6729), .Z(n6727) );
  XOR U6527 ( .A(n6454), .B(n6730), .Z(n6448) );
  IV U6528 ( .A(n6453), .Z(n6730) );
  XNOR U6529 ( .A(n6450), .B(n6639), .Z(n6453) );
  AND U6530 ( .A(n10017), .B(n3166), .Z(n6639) );
  XOR U6531 ( .A(n6731), .B(n6732), .Z(n6450) );
  ANDN U6532 ( .A(n6733), .B(n6734), .Z(n6732) );
  XNOR U6533 ( .A(n6731), .B(n6735), .Z(n6733) );
  XOR U6534 ( .A(n6460), .B(n6736), .Z(n6454) );
  IV U6535 ( .A(n6459), .Z(n6736) );
  XNOR U6536 ( .A(n6456), .B(n6632), .Z(n6459) );
  AND U6537 ( .A(n10387), .B(n2765), .Z(n6632) );
  XOR U6538 ( .A(n6737), .B(n6738), .Z(n6456) );
  ANDN U6539 ( .A(n6739), .B(n6740), .Z(n6738) );
  XNOR U6540 ( .A(n6737), .B(n6741), .Z(n6739) );
  XOR U6541 ( .A(n6466), .B(n6742), .Z(n6460) );
  IV U6542 ( .A(n6465), .Z(n6742) );
  XNOR U6543 ( .A(n6462), .B(n6625), .Z(n6465) );
  AND U6544 ( .A(n10731), .B(n2396), .Z(n6625) );
  XOR U6545 ( .A(n6743), .B(n6744), .Z(n6462) );
  ANDN U6546 ( .A(n6745), .B(n6746), .Z(n6744) );
  XNOR U6547 ( .A(n6743), .B(n6747), .Z(n6745) );
  XOR U6548 ( .A(n6472), .B(n6748), .Z(n6466) );
  IV U6549 ( .A(n6471), .Z(n6748) );
  XNOR U6550 ( .A(n6468), .B(n6618), .Z(n6471) );
  AND U6551 ( .A(n11049), .B(n2053), .Z(n6618) );
  XOR U6552 ( .A(n6749), .B(n6750), .Z(n6468) );
  ANDN U6553 ( .A(n6751), .B(n6752), .Z(n6750) );
  XNOR U6554 ( .A(n6749), .B(n6753), .Z(n6751) );
  XOR U6555 ( .A(n6478), .B(n6754), .Z(n6472) );
  IV U6556 ( .A(n6477), .Z(n6754) );
  XNOR U6557 ( .A(n6474), .B(n6611), .Z(n6477) );
  AND U6558 ( .A(n11341), .B(n1737), .Z(n6611) );
  XOR U6559 ( .A(n6755), .B(n6756), .Z(n6474) );
  ANDN U6560 ( .A(n6757), .B(n6758), .Z(n6756) );
  XNOR U6561 ( .A(n6755), .B(n6759), .Z(n6757) );
  XOR U6562 ( .A(n6484), .B(n6760), .Z(n6478) );
  IV U6563 ( .A(n6483), .Z(n6760) );
  XNOR U6564 ( .A(n6480), .B(n6604), .Z(n6483) );
  AND U6565 ( .A(n11607), .B(n1448), .Z(n6604) );
  XOR U6566 ( .A(n6761), .B(n6762), .Z(n6480) );
  ANDN U6567 ( .A(n6763), .B(n6764), .Z(n6762) );
  XNOR U6568 ( .A(n6761), .B(n6765), .Z(n6763) );
  XOR U6569 ( .A(n6490), .B(n6766), .Z(n6484) );
  IV U6570 ( .A(n6489), .Z(n6766) );
  XNOR U6571 ( .A(n6486), .B(n6597), .Z(n6489) );
  AND U6572 ( .A(n11869), .B(n1185), .Z(n6597) );
  XOR U6573 ( .A(n6767), .B(n6768), .Z(n6486) );
  ANDN U6574 ( .A(n6769), .B(n6770), .Z(n6768) );
  XNOR U6575 ( .A(n6767), .B(n6771), .Z(n6769) );
  XOR U6576 ( .A(n6496), .B(n6772), .Z(n6490) );
  IV U6577 ( .A(n6495), .Z(n6772) );
  XNOR U6578 ( .A(n6492), .B(n6590), .Z(n6495) );
  AND U6579 ( .A(n12128), .B(n948), .Z(n6590) );
  XOR U6580 ( .A(n6773), .B(n6774), .Z(n6492) );
  ANDN U6581 ( .A(n6775), .B(n6776), .Z(n6774) );
  XNOR U6582 ( .A(n6773), .B(n6777), .Z(n6775) );
  XOR U6583 ( .A(n6502), .B(n6778), .Z(n6496) );
  IV U6584 ( .A(n6501), .Z(n6778) );
  XNOR U6585 ( .A(n6498), .B(n6583), .Z(n6501) );
  AND U6586 ( .A(n12387), .B(n736), .Z(n6583) );
  XOR U6587 ( .A(n6779), .B(n6780), .Z(n6498) );
  ANDN U6588 ( .A(n6781), .B(n6782), .Z(n6780) );
  XNOR U6589 ( .A(n6779), .B(n6783), .Z(n6781) );
  XOR U6590 ( .A(n6508), .B(n6784), .Z(n6502) );
  IV U6591 ( .A(n6507), .Z(n6784) );
  XNOR U6592 ( .A(n6504), .B(n6576), .Z(n6507) );
  AND U6593 ( .A(n12644), .B(n552), .Z(n6576) );
  XOR U6594 ( .A(n6785), .B(n6786), .Z(n6504) );
  ANDN U6595 ( .A(n6787), .B(n6788), .Z(n6786) );
  XNOR U6596 ( .A(n6785), .B(n6789), .Z(n6787) );
  XOR U6597 ( .A(n6514), .B(n6790), .Z(n6508) );
  IV U6598 ( .A(n6513), .Z(n6790) );
  XNOR U6599 ( .A(n6510), .B(n6569), .Z(n6513) );
  AND U6600 ( .A(n12880), .B(n395), .Z(n6569) );
  XOR U6601 ( .A(n6791), .B(n6792), .Z(n6510) );
  ANDN U6602 ( .A(n6793), .B(n6794), .Z(n6792) );
  XNOR U6603 ( .A(n6791), .B(n6795), .Z(n6793) );
  XOR U6604 ( .A(n6520), .B(n6796), .Z(n6514) );
  IV U6605 ( .A(n6519), .Z(n6796) );
  XNOR U6606 ( .A(n6516), .B(n6562), .Z(n6519) );
  AND U6607 ( .A(n13070), .B(n264), .Z(n6562) );
  XOR U6608 ( .A(n6797), .B(n6798), .Z(n6516) );
  ANDN U6609 ( .A(n6799), .B(n6800), .Z(n6798) );
  XNOR U6610 ( .A(n6797), .B(n6801), .Z(n6799) );
  XOR U6611 ( .A(n6525), .B(n6802), .Z(n6520) );
  IV U6612 ( .A(n6524), .Z(n6802) );
  XNOR U6613 ( .A(n6521), .B(n6555), .Z(n6524) );
  AND U6614 ( .A(n13207), .B(n159), .Z(n6555) );
  XOR U6615 ( .A(n6803), .B(n6804), .Z(n6521) );
  ANDN U6616 ( .A(n6805), .B(n6806), .Z(n6804) );
  XNOR U6617 ( .A(n6803), .B(n6807), .Z(n6805) );
  XNOR U6618 ( .A(n6531), .B(n6532), .Z(n6525) );
  NANDN U6619 ( .B(n6808), .A(n42), .Z(n6532) );
  XOR U6620 ( .A(n6809), .B(n6810), .Z(n42) );
  XNOR U6621 ( .A(n6528), .B(n6811), .Z(n6531) );
  AND U6622 ( .A(n6527), .B(n80), .Z(n6811) );
  XOR U6623 ( .A(n6812), .B(n6813), .Z(n6528) );
  ANDN U6624 ( .A(n6814), .B(n6815), .Z(n6813) );
  XNOR U6625 ( .A(n6552), .B(n6812), .Z(n6814) );
  XOR U6626 ( .A(n6816), .B(n6539), .Z(n6549) );
  OR U6627 ( .A(n43), .B(n6808), .Z(n6539) );
  XNOR U6628 ( .A(n6809), .B(n6810), .Z(n43) );
  AND U6629 ( .A(n6809), .B(n6817), .Z(n6810) );
  XNOR U6630 ( .A(n6818), .B(n6819), .Z(n6817) );
  ANDN U6631 ( .A(n6819), .B(n6820), .Z(n6818) );
  IV U6632 ( .A(n6533), .Z(n6816) );
  XOR U6633 ( .A(n6821), .B(n6822), .Z(n6533) );
  AND U6634 ( .A(n6823), .B(n6824), .Z(n6822) );
  XOR U6635 ( .A(n6825), .B(n6821), .Z(n6824) );
  XOR U6636 ( .A(n6537), .B(n6545), .Z(n6548) );
  XOR U6637 ( .A(n6826), .B(n6827), .Z(n6537) );
  IV U6638 ( .A(n6828), .Z(n6827) );
  XOR U6639 ( .A(n6829), .B(n6830), .Z(n6545) );
  AND U6640 ( .A(n6829), .B(n6831), .Z(n6830) );
  XOR U6641 ( .A(n6832), .B(n6823), .Z(n6831) );
  XOR U6642 ( .A(n6833), .B(n6553), .Z(n6823) );
  XOR U6643 ( .A(n6560), .B(n6834), .Z(n6553) );
  IV U6644 ( .A(n6558), .Z(n6834) );
  XNOR U6645 ( .A(n6835), .B(n6557), .Z(n6558) );
  OR U6646 ( .A(n6836), .B(n6837), .Z(n6557) );
  NANDN U6647 ( .B(n6541), .A(n159), .Z(n6835) );
  XOR U6648 ( .A(n6567), .B(n6838), .Z(n6560) );
  IV U6649 ( .A(n6566), .Z(n6838) );
  XNOR U6650 ( .A(n6563), .B(n6839), .Z(n6566) );
  XOR U6651 ( .A(n6840), .B(n6841), .Z(n6563) );
  NANDN U6652 ( .B(n6842), .A(n6843), .Z(n6840) );
  XOR U6653 ( .A(n6841), .B(n6844), .Z(n6843) );
  XOR U6654 ( .A(n6574), .B(n6845), .Z(n6567) );
  IV U6655 ( .A(n6573), .Z(n6845) );
  XNOR U6656 ( .A(n6570), .B(n6846), .Z(n6573) );
  XOR U6657 ( .A(n6847), .B(n6848), .Z(n6570) );
  ANDN U6658 ( .A(n6849), .B(n6850), .Z(n6848) );
  XNOR U6659 ( .A(n6847), .B(n6851), .Z(n6849) );
  XOR U6660 ( .A(n6581), .B(n6852), .Z(n6574) );
  IV U6661 ( .A(n6580), .Z(n6852) );
  XNOR U6662 ( .A(n6577), .B(n6853), .Z(n6580) );
  XOR U6663 ( .A(n6854), .B(n6855), .Z(n6577) );
  ANDN U6664 ( .A(n6856), .B(n6857), .Z(n6855) );
  XNOR U6665 ( .A(n6854), .B(n6858), .Z(n6856) );
  XOR U6666 ( .A(n6588), .B(n6859), .Z(n6581) );
  IV U6667 ( .A(n6587), .Z(n6859) );
  XNOR U6668 ( .A(n6584), .B(n6860), .Z(n6587) );
  XOR U6669 ( .A(n6861), .B(n6862), .Z(n6584) );
  ANDN U6670 ( .A(n6863), .B(n6864), .Z(n6862) );
  XNOR U6671 ( .A(n6861), .B(n6865), .Z(n6863) );
  XOR U6672 ( .A(n6595), .B(n6866), .Z(n6588) );
  IV U6673 ( .A(n6594), .Z(n6866) );
  XNOR U6674 ( .A(n6591), .B(n6867), .Z(n6594) );
  XOR U6675 ( .A(n6868), .B(n6869), .Z(n6591) );
  ANDN U6676 ( .A(n6870), .B(n6871), .Z(n6869) );
  XNOR U6677 ( .A(n6868), .B(n6872), .Z(n6870) );
  XOR U6678 ( .A(n6602), .B(n6873), .Z(n6595) );
  IV U6679 ( .A(n6601), .Z(n6873) );
  XNOR U6680 ( .A(n6598), .B(n6874), .Z(n6601) );
  XOR U6681 ( .A(n6875), .B(n6876), .Z(n6598) );
  ANDN U6682 ( .A(n6877), .B(n6878), .Z(n6876) );
  XNOR U6683 ( .A(n6875), .B(n6879), .Z(n6877) );
  XOR U6684 ( .A(n6609), .B(n6880), .Z(n6602) );
  IV U6685 ( .A(n6608), .Z(n6880) );
  XNOR U6686 ( .A(n6605), .B(n6881), .Z(n6608) );
  XOR U6687 ( .A(n6882), .B(n6883), .Z(n6605) );
  ANDN U6688 ( .A(n6884), .B(n6885), .Z(n6883) );
  XNOR U6689 ( .A(n6882), .B(n6886), .Z(n6884) );
  XOR U6690 ( .A(n6616), .B(n6887), .Z(n6609) );
  IV U6691 ( .A(n6615), .Z(n6887) );
  XNOR U6692 ( .A(n6612), .B(n6888), .Z(n6615) );
  XOR U6693 ( .A(n6889), .B(n6890), .Z(n6612) );
  ANDN U6694 ( .A(n6891), .B(n6892), .Z(n6890) );
  XNOR U6695 ( .A(n6889), .B(n6893), .Z(n6891) );
  XOR U6696 ( .A(n6623), .B(n6894), .Z(n6616) );
  IV U6697 ( .A(n6622), .Z(n6894) );
  XNOR U6698 ( .A(n6619), .B(n6895), .Z(n6622) );
  XOR U6699 ( .A(n6896), .B(n6897), .Z(n6619) );
  ANDN U6700 ( .A(n6898), .B(n6899), .Z(n6897) );
  XNOR U6701 ( .A(n6896), .B(n6900), .Z(n6898) );
  XOR U6702 ( .A(n6630), .B(n6901), .Z(n6623) );
  IV U6703 ( .A(n6629), .Z(n6901) );
  XNOR U6704 ( .A(n6626), .B(n6902), .Z(n6629) );
  XOR U6705 ( .A(n6903), .B(n6904), .Z(n6626) );
  ANDN U6706 ( .A(n6905), .B(n6906), .Z(n6904) );
  XNOR U6707 ( .A(n6903), .B(n6907), .Z(n6905) );
  XOR U6708 ( .A(n6637), .B(n6908), .Z(n6630) );
  IV U6709 ( .A(n6636), .Z(n6908) );
  XNOR U6710 ( .A(n6633), .B(n6909), .Z(n6636) );
  XOR U6711 ( .A(n6910), .B(n6911), .Z(n6633) );
  ANDN U6712 ( .A(n6912), .B(n6913), .Z(n6911) );
  XNOR U6713 ( .A(n6910), .B(n6914), .Z(n6912) );
  XOR U6714 ( .A(n6644), .B(n6915), .Z(n6637) );
  IV U6715 ( .A(n6643), .Z(n6915) );
  XNOR U6716 ( .A(n6640), .B(n6916), .Z(n6643) );
  XOR U6717 ( .A(n6917), .B(n6918), .Z(n6640) );
  ANDN U6718 ( .A(n6919), .B(n6920), .Z(n6918) );
  XNOR U6719 ( .A(n6917), .B(n6921), .Z(n6919) );
  XOR U6720 ( .A(n6651), .B(n6922), .Z(n6644) );
  IV U6721 ( .A(n6650), .Z(n6922) );
  XNOR U6722 ( .A(n6647), .B(n6923), .Z(n6650) );
  XOR U6723 ( .A(n6924), .B(n6925), .Z(n6647) );
  ANDN U6724 ( .A(n6926), .B(n6927), .Z(n6925) );
  XNOR U6725 ( .A(n6924), .B(n6928), .Z(n6926) );
  XOR U6726 ( .A(n6658), .B(n6929), .Z(n6651) );
  IV U6727 ( .A(n6657), .Z(n6929) );
  XNOR U6728 ( .A(n6654), .B(n6930), .Z(n6657) );
  XOR U6729 ( .A(n6931), .B(n6932), .Z(n6654) );
  ANDN U6730 ( .A(n6933), .B(n6934), .Z(n6932) );
  XNOR U6731 ( .A(n6931), .B(n6935), .Z(n6933) );
  XOR U6732 ( .A(n6665), .B(n6936), .Z(n6658) );
  IV U6733 ( .A(n6664), .Z(n6936) );
  XNOR U6734 ( .A(n6661), .B(n6937), .Z(n6664) );
  XOR U6735 ( .A(n6938), .B(n6939), .Z(n6661) );
  ANDN U6736 ( .A(n6940), .B(n6941), .Z(n6939) );
  XNOR U6737 ( .A(n6938), .B(n6942), .Z(n6940) );
  XOR U6738 ( .A(n6672), .B(n6943), .Z(n6665) );
  IV U6739 ( .A(n6671), .Z(n6943) );
  XNOR U6740 ( .A(n6668), .B(n6944), .Z(n6671) );
  XOR U6741 ( .A(n6945), .B(n6946), .Z(n6668) );
  ANDN U6742 ( .A(n6947), .B(n6948), .Z(n6946) );
  XNOR U6743 ( .A(n6945), .B(n6949), .Z(n6947) );
  XOR U6744 ( .A(n6679), .B(n6950), .Z(n6672) );
  IV U6745 ( .A(n6678), .Z(n6950) );
  XNOR U6746 ( .A(n6675), .B(n6951), .Z(n6678) );
  XOR U6747 ( .A(n6952), .B(n6953), .Z(n6675) );
  ANDN U6748 ( .A(n6954), .B(n6955), .Z(n6953) );
  XNOR U6749 ( .A(n6952), .B(n6956), .Z(n6954) );
  XOR U6750 ( .A(n6686), .B(n6957), .Z(n6679) );
  IV U6751 ( .A(n6685), .Z(n6957) );
  XNOR U6752 ( .A(n6682), .B(n6958), .Z(n6685) );
  XOR U6753 ( .A(n6959), .B(n6960), .Z(n6682) );
  ANDN U6754 ( .A(n6961), .B(n6962), .Z(n6960) );
  XNOR U6755 ( .A(n6959), .B(n6963), .Z(n6961) );
  XOR U6756 ( .A(n6693), .B(n6964), .Z(n6686) );
  IV U6757 ( .A(n6692), .Z(n6964) );
  XNOR U6758 ( .A(n6689), .B(n6965), .Z(n6692) );
  XOR U6759 ( .A(n6966), .B(n6967), .Z(n6689) );
  ANDN U6760 ( .A(n6968), .B(n6969), .Z(n6967) );
  XNOR U6761 ( .A(n6966), .B(n6970), .Z(n6968) );
  XOR U6762 ( .A(n6699), .B(n6971), .Z(n6693) );
  IV U6763 ( .A(n6698), .Z(n6971) );
  XNOR U6764 ( .A(n6695), .B(n6965), .Z(n6698) );
  AND U6765 ( .A(n7241), .B(n6688), .Z(n6965) );
  XOR U6766 ( .A(n6972), .B(n6973), .Z(n6695) );
  ANDN U6767 ( .A(n6974), .B(n6975), .Z(n6973) );
  XNOR U6768 ( .A(n6972), .B(n6976), .Z(n6974) );
  XOR U6769 ( .A(n6705), .B(n6977), .Z(n6699) );
  IV U6770 ( .A(n6704), .Z(n6977) );
  XNOR U6771 ( .A(n6701), .B(n6958), .Z(n6704) );
  AND U6772 ( .A(n7770), .B(n6118), .Z(n6958) );
  XOR U6773 ( .A(n6978), .B(n6979), .Z(n6701) );
  ANDN U6774 ( .A(n6980), .B(n6981), .Z(n6979) );
  XNOR U6775 ( .A(n6978), .B(n6982), .Z(n6980) );
  XOR U6776 ( .A(n6711), .B(n6983), .Z(n6705) );
  IV U6777 ( .A(n6710), .Z(n6983) );
  XNOR U6778 ( .A(n6707), .B(n6951), .Z(n6710) );
  AND U6779 ( .A(n8272), .B(n5561), .Z(n6951) );
  XOR U6780 ( .A(n6984), .B(n6985), .Z(n6707) );
  ANDN U6781 ( .A(n6986), .B(n6987), .Z(n6985) );
  XNOR U6782 ( .A(n6984), .B(n6988), .Z(n6986) );
  XOR U6783 ( .A(n6717), .B(n6989), .Z(n6711) );
  IV U6784 ( .A(n6716), .Z(n6989) );
  XNOR U6785 ( .A(n6713), .B(n6944), .Z(n6716) );
  AND U6786 ( .A(n8748), .B(n5030), .Z(n6944) );
  XOR U6787 ( .A(n6990), .B(n6991), .Z(n6713) );
  ANDN U6788 ( .A(n6992), .B(n6993), .Z(n6991) );
  XNOR U6789 ( .A(n6990), .B(n6994), .Z(n6992) );
  XOR U6790 ( .A(n6723), .B(n6995), .Z(n6717) );
  IV U6791 ( .A(n6722), .Z(n6995) );
  XNOR U6792 ( .A(n6719), .B(n6937), .Z(n6722) );
  AND U6793 ( .A(n9198), .B(n4525), .Z(n6937) );
  XOR U6794 ( .A(n6996), .B(n6997), .Z(n6719) );
  ANDN U6795 ( .A(n6998), .B(n6999), .Z(n6997) );
  XNOR U6796 ( .A(n6996), .B(n7000), .Z(n6998) );
  XOR U6797 ( .A(n6729), .B(n7001), .Z(n6723) );
  IV U6798 ( .A(n6728), .Z(n7001) );
  XNOR U6799 ( .A(n6725), .B(n6930), .Z(n6728) );
  AND U6800 ( .A(n9621), .B(n4046), .Z(n6930) );
  XOR U6801 ( .A(n7002), .B(n7003), .Z(n6725) );
  ANDN U6802 ( .A(n7004), .B(n7005), .Z(n7003) );
  XNOR U6803 ( .A(n7002), .B(n7006), .Z(n7004) );
  XOR U6804 ( .A(n6735), .B(n7007), .Z(n6729) );
  IV U6805 ( .A(n6734), .Z(n7007) );
  XNOR U6806 ( .A(n6731), .B(n6923), .Z(n6734) );
  AND U6807 ( .A(n10017), .B(n3593), .Z(n6923) );
  XOR U6808 ( .A(n7008), .B(n7009), .Z(n6731) );
  ANDN U6809 ( .A(n7010), .B(n7011), .Z(n7009) );
  XNOR U6810 ( .A(n7008), .B(n7012), .Z(n7010) );
  XOR U6811 ( .A(n6741), .B(n7013), .Z(n6735) );
  IV U6812 ( .A(n6740), .Z(n7013) );
  XNOR U6813 ( .A(n6737), .B(n6916), .Z(n6740) );
  AND U6814 ( .A(n10387), .B(n3166), .Z(n6916) );
  XOR U6815 ( .A(n7014), .B(n7015), .Z(n6737) );
  ANDN U6816 ( .A(n7016), .B(n7017), .Z(n7015) );
  XNOR U6817 ( .A(n7014), .B(n7018), .Z(n7016) );
  XOR U6818 ( .A(n6747), .B(n7019), .Z(n6741) );
  IV U6819 ( .A(n6746), .Z(n7019) );
  XNOR U6820 ( .A(n6743), .B(n6909), .Z(n6746) );
  AND U6821 ( .A(n10731), .B(n2765), .Z(n6909) );
  XOR U6822 ( .A(n7020), .B(n7021), .Z(n6743) );
  ANDN U6823 ( .A(n7022), .B(n7023), .Z(n7021) );
  XNOR U6824 ( .A(n7020), .B(n7024), .Z(n7022) );
  XOR U6825 ( .A(n6753), .B(n7025), .Z(n6747) );
  IV U6826 ( .A(n6752), .Z(n7025) );
  XNOR U6827 ( .A(n6749), .B(n6902), .Z(n6752) );
  AND U6828 ( .A(n11049), .B(n2396), .Z(n6902) );
  XOR U6829 ( .A(n7026), .B(n7027), .Z(n6749) );
  ANDN U6830 ( .A(n7028), .B(n7029), .Z(n7027) );
  XNOR U6831 ( .A(n7026), .B(n7030), .Z(n7028) );
  XOR U6832 ( .A(n6759), .B(n7031), .Z(n6753) );
  IV U6833 ( .A(n6758), .Z(n7031) );
  XNOR U6834 ( .A(n6755), .B(n6895), .Z(n6758) );
  AND U6835 ( .A(n11341), .B(n2053), .Z(n6895) );
  XOR U6836 ( .A(n7032), .B(n7033), .Z(n6755) );
  ANDN U6837 ( .A(n7034), .B(n7035), .Z(n7033) );
  XNOR U6838 ( .A(n7032), .B(n7036), .Z(n7034) );
  XOR U6839 ( .A(n6765), .B(n7037), .Z(n6759) );
  IV U6840 ( .A(n6764), .Z(n7037) );
  XNOR U6841 ( .A(n6761), .B(n6888), .Z(n6764) );
  AND U6842 ( .A(n11607), .B(n1737), .Z(n6888) );
  XOR U6843 ( .A(n7038), .B(n7039), .Z(n6761) );
  ANDN U6844 ( .A(n7040), .B(n7041), .Z(n7039) );
  XNOR U6845 ( .A(n7038), .B(n7042), .Z(n7040) );
  XOR U6846 ( .A(n6771), .B(n7043), .Z(n6765) );
  IV U6847 ( .A(n6770), .Z(n7043) );
  XNOR U6848 ( .A(n6767), .B(n6881), .Z(n6770) );
  AND U6849 ( .A(n11869), .B(n1448), .Z(n6881) );
  XOR U6850 ( .A(n7044), .B(n7045), .Z(n6767) );
  ANDN U6851 ( .A(n7046), .B(n7047), .Z(n7045) );
  XNOR U6852 ( .A(n7044), .B(n7048), .Z(n7046) );
  XOR U6853 ( .A(n6777), .B(n7049), .Z(n6771) );
  IV U6854 ( .A(n6776), .Z(n7049) );
  XNOR U6855 ( .A(n6773), .B(n6874), .Z(n6776) );
  AND U6856 ( .A(n12128), .B(n1185), .Z(n6874) );
  XOR U6857 ( .A(n7050), .B(n7051), .Z(n6773) );
  ANDN U6858 ( .A(n7052), .B(n7053), .Z(n7051) );
  XNOR U6859 ( .A(n7050), .B(n7054), .Z(n7052) );
  XOR U6860 ( .A(n6783), .B(n7055), .Z(n6777) );
  IV U6861 ( .A(n6782), .Z(n7055) );
  XNOR U6862 ( .A(n6779), .B(n6867), .Z(n6782) );
  AND U6863 ( .A(n12387), .B(n948), .Z(n6867) );
  XOR U6864 ( .A(n7056), .B(n7057), .Z(n6779) );
  ANDN U6865 ( .A(n7058), .B(n7059), .Z(n7057) );
  XNOR U6866 ( .A(n7056), .B(n7060), .Z(n7058) );
  XOR U6867 ( .A(n6789), .B(n7061), .Z(n6783) );
  IV U6868 ( .A(n6788), .Z(n7061) );
  XNOR U6869 ( .A(n6785), .B(n6860), .Z(n6788) );
  AND U6870 ( .A(n12644), .B(n736), .Z(n6860) );
  XOR U6871 ( .A(n7062), .B(n7063), .Z(n6785) );
  ANDN U6872 ( .A(n7064), .B(n7065), .Z(n7063) );
  XNOR U6873 ( .A(n7062), .B(n7066), .Z(n7064) );
  XOR U6874 ( .A(n6795), .B(n7067), .Z(n6789) );
  IV U6875 ( .A(n6794), .Z(n7067) );
  XNOR U6876 ( .A(n6791), .B(n6853), .Z(n6794) );
  AND U6877 ( .A(n12880), .B(n552), .Z(n6853) );
  XOR U6878 ( .A(n7068), .B(n7069), .Z(n6791) );
  ANDN U6879 ( .A(n7070), .B(n7071), .Z(n7069) );
  XNOR U6880 ( .A(n7068), .B(n7072), .Z(n7070) );
  XOR U6881 ( .A(n6801), .B(n7073), .Z(n6795) );
  IV U6882 ( .A(n6800), .Z(n7073) );
  XNOR U6883 ( .A(n6797), .B(n6846), .Z(n6800) );
  AND U6884 ( .A(n13070), .B(n395), .Z(n6846) );
  XOR U6885 ( .A(n7074), .B(n7075), .Z(n6797) );
  ANDN U6886 ( .A(n7076), .B(n7077), .Z(n7075) );
  XNOR U6887 ( .A(n7074), .B(n7078), .Z(n7076) );
  XOR U6888 ( .A(n6807), .B(n7079), .Z(n6801) );
  IV U6889 ( .A(n6806), .Z(n7079) );
  XNOR U6890 ( .A(n6803), .B(n6839), .Z(n6806) );
  AND U6891 ( .A(n13207), .B(n264), .Z(n6839) );
  XOR U6892 ( .A(n7080), .B(n7081), .Z(n6803) );
  ANDN U6893 ( .A(n7082), .B(n7083), .Z(n7081) );
  XNOR U6894 ( .A(n7080), .B(n7084), .Z(n7082) );
  XNOR U6895 ( .A(n6815), .B(n6552), .Z(n6807) );
  XNOR U6896 ( .A(n6812), .B(n7085), .Z(n6815) );
  AND U6897 ( .A(n6527), .B(n159), .Z(n7085) );
  XOR U6898 ( .A(n7086), .B(n7087), .Z(n6812) );
  ANDN U6899 ( .A(n7088), .B(n7089), .Z(n7087) );
  XNOR U6900 ( .A(n6836), .B(n7086), .Z(n7088) );
  XOR U6901 ( .A(n7090), .B(n6552), .Z(n6833) );
  NANDN U6902 ( .B(n6808), .A(n80), .Z(n6552) );
  XOR U6903 ( .A(n7091), .B(n7092), .Z(n80) );
  AND U6904 ( .A(n6809), .B(n7093), .Z(n7092) );
  XNOR U6905 ( .A(n7091), .B(n6820), .Z(n7093) );
  XOR U6906 ( .A(n6819), .B(n7091), .Z(n6820) );
  XOR U6907 ( .A(n7094), .B(n7095), .Z(n6819) );
  ANDN U6908 ( .A(n7094), .B(n7096), .Z(n7095) );
  IV U6909 ( .A(n6821), .Z(n7090) );
  XOR U6910 ( .A(n7097), .B(n7098), .Z(n6821) );
  AND U6911 ( .A(n7099), .B(n7100), .Z(n7098) );
  XOR U6912 ( .A(n7101), .B(n7097), .Z(n7100) );
  XOR U6913 ( .A(n6825), .B(n6829), .Z(n6832) );
  XOR U6914 ( .A(n7102), .B(n7103), .Z(n6825) );
  IV U6915 ( .A(n7104), .Z(n7103) );
  XOR U6916 ( .A(n7105), .B(n7106), .Z(n6829) );
  AND U6917 ( .A(n7105), .B(n7107), .Z(n7106) );
  XOR U6918 ( .A(n7108), .B(n7099), .Z(n7107) );
  XOR U6919 ( .A(n7109), .B(n6837), .Z(n7099) );
  XOR U6920 ( .A(n6844), .B(n7110), .Z(n6837) );
  IV U6921 ( .A(n6842), .Z(n7110) );
  XNOR U6922 ( .A(n7111), .B(n6841), .Z(n6842) );
  OR U6923 ( .A(n7112), .B(n7113), .Z(n6841) );
  NANDN U6924 ( .B(n6541), .A(n264), .Z(n7111) );
  XOR U6925 ( .A(n6851), .B(n7114), .Z(n6844) );
  IV U6926 ( .A(n6850), .Z(n7114) );
  XNOR U6927 ( .A(n6847), .B(n7115), .Z(n6850) );
  XOR U6928 ( .A(n7116), .B(n7117), .Z(n6847) );
  NANDN U6929 ( .B(n7118), .A(n7119), .Z(n7116) );
  XOR U6930 ( .A(n7117), .B(n7120), .Z(n7119) );
  XOR U6931 ( .A(n6858), .B(n7121), .Z(n6851) );
  IV U6932 ( .A(n6857), .Z(n7121) );
  XNOR U6933 ( .A(n6854), .B(n7122), .Z(n6857) );
  XOR U6934 ( .A(n7123), .B(n7124), .Z(n6854) );
  ANDN U6935 ( .A(n7125), .B(n7126), .Z(n7124) );
  XNOR U6936 ( .A(n7123), .B(n7127), .Z(n7125) );
  XOR U6937 ( .A(n6865), .B(n7128), .Z(n6858) );
  IV U6938 ( .A(n6864), .Z(n7128) );
  XNOR U6939 ( .A(n6861), .B(n7129), .Z(n6864) );
  XOR U6940 ( .A(n7130), .B(n7131), .Z(n6861) );
  ANDN U6941 ( .A(n7132), .B(n7133), .Z(n7131) );
  XNOR U6942 ( .A(n7130), .B(n7134), .Z(n7132) );
  XOR U6943 ( .A(n6872), .B(n7135), .Z(n6865) );
  IV U6944 ( .A(n6871), .Z(n7135) );
  XNOR U6945 ( .A(n6868), .B(n7136), .Z(n6871) );
  XOR U6946 ( .A(n7137), .B(n7138), .Z(n6868) );
  ANDN U6947 ( .A(n7139), .B(n7140), .Z(n7138) );
  XNOR U6948 ( .A(n7137), .B(n7141), .Z(n7139) );
  XOR U6949 ( .A(n6879), .B(n7142), .Z(n6872) );
  IV U6950 ( .A(n6878), .Z(n7142) );
  XNOR U6951 ( .A(n6875), .B(n7143), .Z(n6878) );
  XOR U6952 ( .A(n7144), .B(n7145), .Z(n6875) );
  ANDN U6953 ( .A(n7146), .B(n7147), .Z(n7145) );
  XNOR U6954 ( .A(n7144), .B(n7148), .Z(n7146) );
  XOR U6955 ( .A(n6886), .B(n7149), .Z(n6879) );
  IV U6956 ( .A(n6885), .Z(n7149) );
  XNOR U6957 ( .A(n6882), .B(n7150), .Z(n6885) );
  XOR U6958 ( .A(n7151), .B(n7152), .Z(n6882) );
  ANDN U6959 ( .A(n7153), .B(n7154), .Z(n7152) );
  XNOR U6960 ( .A(n7151), .B(n7155), .Z(n7153) );
  XOR U6961 ( .A(n6893), .B(n7156), .Z(n6886) );
  IV U6962 ( .A(n6892), .Z(n7156) );
  XNOR U6963 ( .A(n6889), .B(n7157), .Z(n6892) );
  XOR U6964 ( .A(n7158), .B(n7159), .Z(n6889) );
  ANDN U6965 ( .A(n7160), .B(n7161), .Z(n7159) );
  XNOR U6966 ( .A(n7158), .B(n7162), .Z(n7160) );
  XOR U6967 ( .A(n6900), .B(n7163), .Z(n6893) );
  IV U6968 ( .A(n6899), .Z(n7163) );
  XNOR U6969 ( .A(n6896), .B(n7164), .Z(n6899) );
  XOR U6970 ( .A(n7165), .B(n7166), .Z(n6896) );
  ANDN U6971 ( .A(n7167), .B(n7168), .Z(n7166) );
  XNOR U6972 ( .A(n7165), .B(n7169), .Z(n7167) );
  XOR U6973 ( .A(n6907), .B(n7170), .Z(n6900) );
  IV U6974 ( .A(n6906), .Z(n7170) );
  XNOR U6975 ( .A(n6903), .B(n7171), .Z(n6906) );
  XOR U6976 ( .A(n7172), .B(n7173), .Z(n6903) );
  ANDN U6977 ( .A(n7174), .B(n7175), .Z(n7173) );
  XNOR U6978 ( .A(n7172), .B(n7176), .Z(n7174) );
  XOR U6979 ( .A(n6914), .B(n7177), .Z(n6907) );
  IV U6980 ( .A(n6913), .Z(n7177) );
  XNOR U6981 ( .A(n6910), .B(n7178), .Z(n6913) );
  XOR U6982 ( .A(n7179), .B(n7180), .Z(n6910) );
  ANDN U6983 ( .A(n7181), .B(n7182), .Z(n7180) );
  XNOR U6984 ( .A(n7179), .B(n7183), .Z(n7181) );
  XOR U6985 ( .A(n6921), .B(n7184), .Z(n6914) );
  IV U6986 ( .A(n6920), .Z(n7184) );
  XNOR U6987 ( .A(n6917), .B(n7185), .Z(n6920) );
  XOR U6988 ( .A(n7186), .B(n7187), .Z(n6917) );
  ANDN U6989 ( .A(n7188), .B(n7189), .Z(n7187) );
  XNOR U6990 ( .A(n7186), .B(n7190), .Z(n7188) );
  XOR U6991 ( .A(n6928), .B(n7191), .Z(n6921) );
  IV U6992 ( .A(n6927), .Z(n7191) );
  XNOR U6993 ( .A(n6924), .B(n7192), .Z(n6927) );
  XOR U6994 ( .A(n7193), .B(n7194), .Z(n6924) );
  ANDN U6995 ( .A(n7195), .B(n7196), .Z(n7194) );
  XNOR U6996 ( .A(n7193), .B(n7197), .Z(n7195) );
  XOR U6997 ( .A(n6935), .B(n7198), .Z(n6928) );
  IV U6998 ( .A(n6934), .Z(n7198) );
  XNOR U6999 ( .A(n6931), .B(n7199), .Z(n6934) );
  XOR U7000 ( .A(n7200), .B(n7201), .Z(n6931) );
  ANDN U7001 ( .A(n7202), .B(n7203), .Z(n7201) );
  XNOR U7002 ( .A(n7200), .B(n7204), .Z(n7202) );
  XOR U7003 ( .A(n6942), .B(n7205), .Z(n6935) );
  IV U7004 ( .A(n6941), .Z(n7205) );
  XNOR U7005 ( .A(n6938), .B(n7206), .Z(n6941) );
  XOR U7006 ( .A(n7207), .B(n7208), .Z(n6938) );
  ANDN U7007 ( .A(n7209), .B(n7210), .Z(n7208) );
  XNOR U7008 ( .A(n7207), .B(n7211), .Z(n7209) );
  XOR U7009 ( .A(n6949), .B(n7212), .Z(n6942) );
  IV U7010 ( .A(n6948), .Z(n7212) );
  XNOR U7011 ( .A(n6945), .B(n7213), .Z(n6948) );
  XOR U7012 ( .A(n7214), .B(n7215), .Z(n6945) );
  ANDN U7013 ( .A(n7216), .B(n7217), .Z(n7215) );
  XNOR U7014 ( .A(n7214), .B(n7218), .Z(n7216) );
  XOR U7015 ( .A(n6956), .B(n7219), .Z(n6949) );
  IV U7016 ( .A(n6955), .Z(n7219) );
  XNOR U7017 ( .A(n6952), .B(n7220), .Z(n6955) );
  XOR U7018 ( .A(n7221), .B(n7222), .Z(n6952) );
  ANDN U7019 ( .A(n7223), .B(n7224), .Z(n7222) );
  XNOR U7020 ( .A(n7221), .B(n7225), .Z(n7223) );
  XOR U7021 ( .A(n6963), .B(n7226), .Z(n6956) );
  IV U7022 ( .A(n6962), .Z(n7226) );
  XNOR U7023 ( .A(n6959), .B(n7227), .Z(n6962) );
  XOR U7024 ( .A(n7228), .B(n7229), .Z(n6959) );
  ANDN U7025 ( .A(n7230), .B(n7231), .Z(n7229) );
  XNOR U7026 ( .A(n7228), .B(n7232), .Z(n7230) );
  XOR U7027 ( .A(n6970), .B(n7233), .Z(n6963) );
  IV U7028 ( .A(n6969), .Z(n7233) );
  XNOR U7029 ( .A(n6966), .B(n7234), .Z(n6969) );
  XOR U7030 ( .A(n7235), .B(n7236), .Z(n6966) );
  ANDN U7031 ( .A(n7237), .B(n7238), .Z(n7236) );
  XNOR U7032 ( .A(n7235), .B(n7239), .Z(n7237) );
  XOR U7033 ( .A(n6976), .B(n7240), .Z(n6970) );
  IV U7034 ( .A(n6975), .Z(n7240) );
  XNOR U7035 ( .A(n6972), .B(n7241), .Z(n6975) );
  XOR U7036 ( .A(n7242), .B(n7243), .Z(n6972) );
  ANDN U7037 ( .A(n7244), .B(n7245), .Z(n7243) );
  XNOR U7038 ( .A(n7242), .B(n7246), .Z(n7244) );
  XOR U7039 ( .A(n6982), .B(n7247), .Z(n6976) );
  IV U7040 ( .A(n6981), .Z(n7247) );
  XNOR U7041 ( .A(n6978), .B(n7234), .Z(n6981) );
  AND U7042 ( .A(n7770), .B(n6688), .Z(n7234) );
  XOR U7043 ( .A(n7248), .B(n7249), .Z(n6978) );
  ANDN U7044 ( .A(n7250), .B(n7251), .Z(n7249) );
  XNOR U7045 ( .A(n7248), .B(n7252), .Z(n7250) );
  XOR U7046 ( .A(n6988), .B(n7253), .Z(n6982) );
  IV U7047 ( .A(n6987), .Z(n7253) );
  XNOR U7048 ( .A(n6984), .B(n7227), .Z(n6987) );
  AND U7049 ( .A(n8272), .B(n6118), .Z(n7227) );
  XOR U7050 ( .A(n7254), .B(n7255), .Z(n6984) );
  ANDN U7051 ( .A(n7256), .B(n7257), .Z(n7255) );
  XNOR U7052 ( .A(n7254), .B(n7258), .Z(n7256) );
  XOR U7053 ( .A(n6994), .B(n7259), .Z(n6988) );
  IV U7054 ( .A(n6993), .Z(n7259) );
  XNOR U7055 ( .A(n6990), .B(n7220), .Z(n6993) );
  AND U7056 ( .A(n8748), .B(n5561), .Z(n7220) );
  XOR U7057 ( .A(n7260), .B(n7261), .Z(n6990) );
  ANDN U7058 ( .A(n7262), .B(n7263), .Z(n7261) );
  XNOR U7059 ( .A(n7260), .B(n7264), .Z(n7262) );
  XOR U7060 ( .A(n7000), .B(n7265), .Z(n6994) );
  IV U7061 ( .A(n6999), .Z(n7265) );
  XNOR U7062 ( .A(n6996), .B(n7213), .Z(n6999) );
  AND U7063 ( .A(n9198), .B(n5030), .Z(n7213) );
  XOR U7064 ( .A(n7266), .B(n7267), .Z(n6996) );
  ANDN U7065 ( .A(n7268), .B(n7269), .Z(n7267) );
  XNOR U7066 ( .A(n7266), .B(n7270), .Z(n7268) );
  XOR U7067 ( .A(n7006), .B(n7271), .Z(n7000) );
  IV U7068 ( .A(n7005), .Z(n7271) );
  XNOR U7069 ( .A(n7002), .B(n7206), .Z(n7005) );
  AND U7070 ( .A(n9621), .B(n4525), .Z(n7206) );
  XOR U7071 ( .A(n7272), .B(n7273), .Z(n7002) );
  ANDN U7072 ( .A(n7274), .B(n7275), .Z(n7273) );
  XNOR U7073 ( .A(n7272), .B(n7276), .Z(n7274) );
  XOR U7074 ( .A(n7012), .B(n7277), .Z(n7006) );
  IV U7075 ( .A(n7011), .Z(n7277) );
  XNOR U7076 ( .A(n7008), .B(n7199), .Z(n7011) );
  AND U7077 ( .A(n10017), .B(n4046), .Z(n7199) );
  XOR U7078 ( .A(n7278), .B(n7279), .Z(n7008) );
  ANDN U7079 ( .A(n7280), .B(n7281), .Z(n7279) );
  XNOR U7080 ( .A(n7278), .B(n7282), .Z(n7280) );
  XOR U7081 ( .A(n7018), .B(n7283), .Z(n7012) );
  IV U7082 ( .A(n7017), .Z(n7283) );
  XNOR U7083 ( .A(n7014), .B(n7192), .Z(n7017) );
  AND U7084 ( .A(n10387), .B(n3593), .Z(n7192) );
  XOR U7085 ( .A(n7284), .B(n7285), .Z(n7014) );
  ANDN U7086 ( .A(n7286), .B(n7287), .Z(n7285) );
  XNOR U7087 ( .A(n7284), .B(n7288), .Z(n7286) );
  XOR U7088 ( .A(n7024), .B(n7289), .Z(n7018) );
  IV U7089 ( .A(n7023), .Z(n7289) );
  XNOR U7090 ( .A(n7020), .B(n7185), .Z(n7023) );
  AND U7091 ( .A(n10731), .B(n3166), .Z(n7185) );
  XOR U7092 ( .A(n7290), .B(n7291), .Z(n7020) );
  ANDN U7093 ( .A(n7292), .B(n7293), .Z(n7291) );
  XNOR U7094 ( .A(n7290), .B(n7294), .Z(n7292) );
  XOR U7095 ( .A(n7030), .B(n7295), .Z(n7024) );
  IV U7096 ( .A(n7029), .Z(n7295) );
  XNOR U7097 ( .A(n7026), .B(n7178), .Z(n7029) );
  AND U7098 ( .A(n11049), .B(n2765), .Z(n7178) );
  XOR U7099 ( .A(n7296), .B(n7297), .Z(n7026) );
  ANDN U7100 ( .A(n7298), .B(n7299), .Z(n7297) );
  XNOR U7101 ( .A(n7296), .B(n7300), .Z(n7298) );
  XOR U7102 ( .A(n7036), .B(n7301), .Z(n7030) );
  IV U7103 ( .A(n7035), .Z(n7301) );
  XNOR U7104 ( .A(n7032), .B(n7171), .Z(n7035) );
  AND U7105 ( .A(n11341), .B(n2396), .Z(n7171) );
  XOR U7106 ( .A(n7302), .B(n7303), .Z(n7032) );
  ANDN U7107 ( .A(n7304), .B(n7305), .Z(n7303) );
  XNOR U7108 ( .A(n7302), .B(n7306), .Z(n7304) );
  XOR U7109 ( .A(n7042), .B(n7307), .Z(n7036) );
  IV U7110 ( .A(n7041), .Z(n7307) );
  XNOR U7111 ( .A(n7038), .B(n7164), .Z(n7041) );
  AND U7112 ( .A(n11607), .B(n2053), .Z(n7164) );
  XOR U7113 ( .A(n7308), .B(n7309), .Z(n7038) );
  ANDN U7114 ( .A(n7310), .B(n7311), .Z(n7309) );
  XNOR U7115 ( .A(n7308), .B(n7312), .Z(n7310) );
  XOR U7116 ( .A(n7048), .B(n7313), .Z(n7042) );
  IV U7117 ( .A(n7047), .Z(n7313) );
  XNOR U7118 ( .A(n7044), .B(n7157), .Z(n7047) );
  AND U7119 ( .A(n11869), .B(n1737), .Z(n7157) );
  XOR U7120 ( .A(n7314), .B(n7315), .Z(n7044) );
  ANDN U7121 ( .A(n7316), .B(n7317), .Z(n7315) );
  XNOR U7122 ( .A(n7314), .B(n7318), .Z(n7316) );
  XOR U7123 ( .A(n7054), .B(n7319), .Z(n7048) );
  IV U7124 ( .A(n7053), .Z(n7319) );
  XNOR U7125 ( .A(n7050), .B(n7150), .Z(n7053) );
  AND U7126 ( .A(n12128), .B(n1448), .Z(n7150) );
  XOR U7127 ( .A(n7320), .B(n7321), .Z(n7050) );
  ANDN U7128 ( .A(n7322), .B(n7323), .Z(n7321) );
  XNOR U7129 ( .A(n7320), .B(n7324), .Z(n7322) );
  XOR U7130 ( .A(n7060), .B(n7325), .Z(n7054) );
  IV U7131 ( .A(n7059), .Z(n7325) );
  XNOR U7132 ( .A(n7056), .B(n7143), .Z(n7059) );
  AND U7133 ( .A(n12387), .B(n1185), .Z(n7143) );
  XOR U7134 ( .A(n7326), .B(n7327), .Z(n7056) );
  ANDN U7135 ( .A(n7328), .B(n7329), .Z(n7327) );
  XNOR U7136 ( .A(n7326), .B(n7330), .Z(n7328) );
  XOR U7137 ( .A(n7066), .B(n7331), .Z(n7060) );
  IV U7138 ( .A(n7065), .Z(n7331) );
  XNOR U7139 ( .A(n7062), .B(n7136), .Z(n7065) );
  AND U7140 ( .A(n12644), .B(n948), .Z(n7136) );
  XOR U7141 ( .A(n7332), .B(n7333), .Z(n7062) );
  ANDN U7142 ( .A(n7334), .B(n7335), .Z(n7333) );
  XNOR U7143 ( .A(n7332), .B(n7336), .Z(n7334) );
  XOR U7144 ( .A(n7072), .B(n7337), .Z(n7066) );
  IV U7145 ( .A(n7071), .Z(n7337) );
  XNOR U7146 ( .A(n7068), .B(n7129), .Z(n7071) );
  AND U7147 ( .A(n12880), .B(n736), .Z(n7129) );
  XOR U7148 ( .A(n7338), .B(n7339), .Z(n7068) );
  ANDN U7149 ( .A(n7340), .B(n7341), .Z(n7339) );
  XNOR U7150 ( .A(n7338), .B(n7342), .Z(n7340) );
  XOR U7151 ( .A(n7078), .B(n7343), .Z(n7072) );
  IV U7152 ( .A(n7077), .Z(n7343) );
  XNOR U7153 ( .A(n7074), .B(n7122), .Z(n7077) );
  AND U7154 ( .A(n13070), .B(n552), .Z(n7122) );
  XOR U7155 ( .A(n7344), .B(n7345), .Z(n7074) );
  ANDN U7156 ( .A(n7346), .B(n7347), .Z(n7345) );
  XNOR U7157 ( .A(n7344), .B(n7348), .Z(n7346) );
  XOR U7158 ( .A(n7084), .B(n7349), .Z(n7078) );
  IV U7159 ( .A(n7083), .Z(n7349) );
  XNOR U7160 ( .A(n7080), .B(n7115), .Z(n7083) );
  AND U7161 ( .A(n13207), .B(n395), .Z(n7115) );
  XOR U7162 ( .A(n7350), .B(n7351), .Z(n7080) );
  ANDN U7163 ( .A(n7352), .B(n7353), .Z(n7351) );
  XNOR U7164 ( .A(n7350), .B(n7354), .Z(n7352) );
  XNOR U7165 ( .A(n7089), .B(n6836), .Z(n7084) );
  XNOR U7166 ( .A(n7086), .B(n7355), .Z(n7089) );
  AND U7167 ( .A(n6527), .B(n264), .Z(n7355) );
  XOR U7168 ( .A(n7356), .B(n7357), .Z(n7086) );
  ANDN U7169 ( .A(n7358), .B(n7359), .Z(n7357) );
  XNOR U7170 ( .A(n7112), .B(n7356), .Z(n7358) );
  XOR U7171 ( .A(n7360), .B(n6836), .Z(n7109) );
  NANDN U7172 ( .B(n6808), .A(n159), .Z(n6836) );
  XOR U7173 ( .A(n7361), .B(n7362), .Z(n159) );
  AND U7174 ( .A(n6809), .B(n7363), .Z(n7362) );
  XNOR U7175 ( .A(n7361), .B(n7096), .Z(n7363) );
  XOR U7176 ( .A(n7094), .B(n7361), .Z(n7096) );
  XOR U7177 ( .A(n7364), .B(n7365), .Z(n7094) );
  ANDN U7178 ( .A(n7364), .B(n7366), .Z(n7365) );
  XOR U7179 ( .A(n7367), .B(n7368), .Z(n7361) );
  IV U7180 ( .A(n7097), .Z(n7360) );
  XOR U7181 ( .A(n7369), .B(n7370), .Z(n7097) );
  AND U7182 ( .A(n7371), .B(n7372), .Z(n7370) );
  XOR U7183 ( .A(n7373), .B(n7369), .Z(n7372) );
  XOR U7184 ( .A(n7101), .B(n7105), .Z(n7108) );
  XOR U7185 ( .A(n7374), .B(n7375), .Z(n7101) );
  IV U7186 ( .A(n7376), .Z(n7375) );
  XOR U7187 ( .A(n7377), .B(n7378), .Z(n7105) );
  AND U7188 ( .A(n7377), .B(n7379), .Z(n7378) );
  XOR U7189 ( .A(n7380), .B(n7371), .Z(n7379) );
  XOR U7190 ( .A(n7381), .B(n7113), .Z(n7371) );
  XOR U7191 ( .A(n7120), .B(n7382), .Z(n7113) );
  IV U7192 ( .A(n7118), .Z(n7382) );
  XNOR U7193 ( .A(n7383), .B(n7117), .Z(n7118) );
  OR U7194 ( .A(n7384), .B(n7385), .Z(n7117) );
  NANDN U7195 ( .B(n6541), .A(n395), .Z(n7383) );
  XOR U7196 ( .A(n7127), .B(n7386), .Z(n7120) );
  IV U7197 ( .A(n7126), .Z(n7386) );
  XNOR U7198 ( .A(n7123), .B(n7387), .Z(n7126) );
  XOR U7199 ( .A(n7388), .B(n7389), .Z(n7123) );
  NANDN U7200 ( .B(n7390), .A(n7391), .Z(n7388) );
  XOR U7201 ( .A(n7389), .B(n7392), .Z(n7391) );
  XOR U7202 ( .A(n7134), .B(n7393), .Z(n7127) );
  IV U7203 ( .A(n7133), .Z(n7393) );
  XNOR U7204 ( .A(n7130), .B(n7394), .Z(n7133) );
  XOR U7205 ( .A(n7395), .B(n7396), .Z(n7130) );
  ANDN U7206 ( .A(n7397), .B(n7398), .Z(n7396) );
  XNOR U7207 ( .A(n7395), .B(n7399), .Z(n7397) );
  XOR U7208 ( .A(n7141), .B(n7400), .Z(n7134) );
  IV U7209 ( .A(n7140), .Z(n7400) );
  XNOR U7210 ( .A(n7137), .B(n7401), .Z(n7140) );
  XOR U7211 ( .A(n7402), .B(n7403), .Z(n7137) );
  ANDN U7212 ( .A(n7404), .B(n7405), .Z(n7403) );
  XNOR U7213 ( .A(n7402), .B(n7406), .Z(n7404) );
  XOR U7214 ( .A(n7148), .B(n7407), .Z(n7141) );
  IV U7215 ( .A(n7147), .Z(n7407) );
  XNOR U7216 ( .A(n7144), .B(n7408), .Z(n7147) );
  XOR U7217 ( .A(n7409), .B(n7410), .Z(n7144) );
  ANDN U7218 ( .A(n7411), .B(n7412), .Z(n7410) );
  XNOR U7219 ( .A(n7409), .B(n7413), .Z(n7411) );
  XOR U7220 ( .A(n7155), .B(n7414), .Z(n7148) );
  IV U7221 ( .A(n7154), .Z(n7414) );
  XNOR U7222 ( .A(n7151), .B(n7415), .Z(n7154) );
  XOR U7223 ( .A(n7416), .B(n7417), .Z(n7151) );
  ANDN U7224 ( .A(n7418), .B(n7419), .Z(n7417) );
  XNOR U7225 ( .A(n7416), .B(n7420), .Z(n7418) );
  XOR U7226 ( .A(n7162), .B(n7421), .Z(n7155) );
  IV U7227 ( .A(n7161), .Z(n7421) );
  XNOR U7228 ( .A(n7158), .B(n7422), .Z(n7161) );
  XOR U7229 ( .A(n7423), .B(n7424), .Z(n7158) );
  ANDN U7230 ( .A(n7425), .B(n7426), .Z(n7424) );
  XNOR U7231 ( .A(n7423), .B(n7427), .Z(n7425) );
  XOR U7232 ( .A(n7169), .B(n7428), .Z(n7162) );
  IV U7233 ( .A(n7168), .Z(n7428) );
  XNOR U7234 ( .A(n7165), .B(n7429), .Z(n7168) );
  XOR U7235 ( .A(n7430), .B(n7431), .Z(n7165) );
  ANDN U7236 ( .A(n7432), .B(n7433), .Z(n7431) );
  XNOR U7237 ( .A(n7430), .B(n7434), .Z(n7432) );
  XOR U7238 ( .A(n7176), .B(n7435), .Z(n7169) );
  IV U7239 ( .A(n7175), .Z(n7435) );
  XNOR U7240 ( .A(n7172), .B(n7436), .Z(n7175) );
  XOR U7241 ( .A(n7437), .B(n7438), .Z(n7172) );
  ANDN U7242 ( .A(n7439), .B(n7440), .Z(n7438) );
  XNOR U7243 ( .A(n7437), .B(n7441), .Z(n7439) );
  XOR U7244 ( .A(n7183), .B(n7442), .Z(n7176) );
  IV U7245 ( .A(n7182), .Z(n7442) );
  XNOR U7246 ( .A(n7179), .B(n7443), .Z(n7182) );
  XOR U7247 ( .A(n7444), .B(n7445), .Z(n7179) );
  ANDN U7248 ( .A(n7446), .B(n7447), .Z(n7445) );
  XNOR U7249 ( .A(n7444), .B(n7448), .Z(n7446) );
  XOR U7250 ( .A(n7190), .B(n7449), .Z(n7183) );
  IV U7251 ( .A(n7189), .Z(n7449) );
  XNOR U7252 ( .A(n7186), .B(n7450), .Z(n7189) );
  XOR U7253 ( .A(n7451), .B(n7452), .Z(n7186) );
  ANDN U7254 ( .A(n7453), .B(n7454), .Z(n7452) );
  XNOR U7255 ( .A(n7451), .B(n7455), .Z(n7453) );
  XOR U7256 ( .A(n7197), .B(n7456), .Z(n7190) );
  IV U7257 ( .A(n7196), .Z(n7456) );
  XNOR U7258 ( .A(n7193), .B(n7457), .Z(n7196) );
  XOR U7259 ( .A(n7458), .B(n7459), .Z(n7193) );
  ANDN U7260 ( .A(n7460), .B(n7461), .Z(n7459) );
  XNOR U7261 ( .A(n7458), .B(n7462), .Z(n7460) );
  XOR U7262 ( .A(n7204), .B(n7463), .Z(n7197) );
  IV U7263 ( .A(n7203), .Z(n7463) );
  XNOR U7264 ( .A(n7200), .B(n7464), .Z(n7203) );
  XOR U7265 ( .A(n7465), .B(n7466), .Z(n7200) );
  ANDN U7266 ( .A(n7467), .B(n7468), .Z(n7466) );
  XNOR U7267 ( .A(n7465), .B(n7469), .Z(n7467) );
  XOR U7268 ( .A(n7211), .B(n7470), .Z(n7204) );
  IV U7269 ( .A(n7210), .Z(n7470) );
  XNOR U7270 ( .A(n7207), .B(n7471), .Z(n7210) );
  XOR U7271 ( .A(n7472), .B(n7473), .Z(n7207) );
  ANDN U7272 ( .A(n7474), .B(n7475), .Z(n7473) );
  XNOR U7273 ( .A(n7472), .B(n7476), .Z(n7474) );
  XOR U7274 ( .A(n7218), .B(n7477), .Z(n7211) );
  IV U7275 ( .A(n7217), .Z(n7477) );
  XNOR U7276 ( .A(n7214), .B(n7478), .Z(n7217) );
  XOR U7277 ( .A(n7479), .B(n7480), .Z(n7214) );
  ANDN U7278 ( .A(n7481), .B(n7482), .Z(n7480) );
  XNOR U7279 ( .A(n7479), .B(n7483), .Z(n7481) );
  XOR U7280 ( .A(n7225), .B(n7484), .Z(n7218) );
  IV U7281 ( .A(n7224), .Z(n7484) );
  XNOR U7282 ( .A(n7221), .B(n7485), .Z(n7224) );
  XOR U7283 ( .A(n7486), .B(n7487), .Z(n7221) );
  ANDN U7284 ( .A(n7488), .B(n7489), .Z(n7487) );
  XNOR U7285 ( .A(n7486), .B(n7490), .Z(n7488) );
  XOR U7286 ( .A(n7232), .B(n7491), .Z(n7225) );
  IV U7287 ( .A(n7231), .Z(n7491) );
  XNOR U7288 ( .A(n7228), .B(n7492), .Z(n7231) );
  XOR U7289 ( .A(n7493), .B(n7494), .Z(n7228) );
  ANDN U7290 ( .A(n7495), .B(n7496), .Z(n7494) );
  XNOR U7291 ( .A(n7493), .B(n7497), .Z(n7495) );
  XOR U7292 ( .A(n7239), .B(n7498), .Z(n7232) );
  IV U7293 ( .A(n7238), .Z(n7498) );
  XNOR U7294 ( .A(n7235), .B(n7499), .Z(n7238) );
  XOR U7295 ( .A(n7500), .B(n7501), .Z(n7235) );
  ANDN U7296 ( .A(n7502), .B(n7503), .Z(n7501) );
  XNOR U7297 ( .A(n7500), .B(n7504), .Z(n7502) );
  XOR U7298 ( .A(n7246), .B(n7505), .Z(n7239) );
  IV U7299 ( .A(n7245), .Z(n7505) );
  XNOR U7300 ( .A(n7242), .B(n7506), .Z(n7245) );
  XOR U7301 ( .A(n7507), .B(n7508), .Z(n7242) );
  ANDN U7302 ( .A(n7509), .B(n7510), .Z(n7508) );
  XNOR U7303 ( .A(n7507), .B(n7511), .Z(n7509) );
  XOR U7304 ( .A(n7252), .B(n7512), .Z(n7246) );
  IV U7305 ( .A(n7251), .Z(n7512) );
  XNOR U7306 ( .A(n7248), .B(n7506), .Z(n7251) );
  AND U7307 ( .A(n7770), .B(n7241), .Z(n7506) );
  XOR U7308 ( .A(n7513), .B(n7514), .Z(n7248) );
  ANDN U7309 ( .A(n7515), .B(n7516), .Z(n7514) );
  XNOR U7310 ( .A(n7513), .B(n7517), .Z(n7515) );
  XOR U7311 ( .A(n7258), .B(n7518), .Z(n7252) );
  IV U7312 ( .A(n7257), .Z(n7518) );
  XNOR U7313 ( .A(n7254), .B(n7499), .Z(n7257) );
  AND U7314 ( .A(n8272), .B(n6688), .Z(n7499) );
  XOR U7315 ( .A(n7519), .B(n7520), .Z(n7254) );
  ANDN U7316 ( .A(n7521), .B(n7522), .Z(n7520) );
  XNOR U7317 ( .A(n7519), .B(n7523), .Z(n7521) );
  XOR U7318 ( .A(n7264), .B(n7524), .Z(n7258) );
  IV U7319 ( .A(n7263), .Z(n7524) );
  XNOR U7320 ( .A(n7260), .B(n7492), .Z(n7263) );
  AND U7321 ( .A(n8748), .B(n6118), .Z(n7492) );
  XOR U7322 ( .A(n7525), .B(n7526), .Z(n7260) );
  ANDN U7323 ( .A(n7527), .B(n7528), .Z(n7526) );
  XNOR U7324 ( .A(n7525), .B(n7529), .Z(n7527) );
  XOR U7325 ( .A(n7270), .B(n7530), .Z(n7264) );
  IV U7326 ( .A(n7269), .Z(n7530) );
  XNOR U7327 ( .A(n7266), .B(n7485), .Z(n7269) );
  AND U7328 ( .A(n9198), .B(n5561), .Z(n7485) );
  XOR U7329 ( .A(n7531), .B(n7532), .Z(n7266) );
  ANDN U7330 ( .A(n7533), .B(n7534), .Z(n7532) );
  XNOR U7331 ( .A(n7531), .B(n7535), .Z(n7533) );
  XOR U7332 ( .A(n7276), .B(n7536), .Z(n7270) );
  IV U7333 ( .A(n7275), .Z(n7536) );
  XNOR U7334 ( .A(n7272), .B(n7478), .Z(n7275) );
  AND U7335 ( .A(n9621), .B(n5030), .Z(n7478) );
  XOR U7336 ( .A(n7537), .B(n7538), .Z(n7272) );
  ANDN U7337 ( .A(n7539), .B(n7540), .Z(n7538) );
  XNOR U7338 ( .A(n7537), .B(n7541), .Z(n7539) );
  XOR U7339 ( .A(n7282), .B(n7542), .Z(n7276) );
  IV U7340 ( .A(n7281), .Z(n7542) );
  XNOR U7341 ( .A(n7278), .B(n7471), .Z(n7281) );
  AND U7342 ( .A(n10017), .B(n4525), .Z(n7471) );
  XOR U7343 ( .A(n7543), .B(n7544), .Z(n7278) );
  ANDN U7344 ( .A(n7545), .B(n7546), .Z(n7544) );
  XNOR U7345 ( .A(n7543), .B(n7547), .Z(n7545) );
  XOR U7346 ( .A(n7288), .B(n7548), .Z(n7282) );
  IV U7347 ( .A(n7287), .Z(n7548) );
  XNOR U7348 ( .A(n7284), .B(n7464), .Z(n7287) );
  AND U7349 ( .A(n10387), .B(n4046), .Z(n7464) );
  XOR U7350 ( .A(n7549), .B(n7550), .Z(n7284) );
  ANDN U7351 ( .A(n7551), .B(n7552), .Z(n7550) );
  XNOR U7352 ( .A(n7549), .B(n7553), .Z(n7551) );
  XOR U7353 ( .A(n7294), .B(n7554), .Z(n7288) );
  IV U7354 ( .A(n7293), .Z(n7554) );
  XNOR U7355 ( .A(n7290), .B(n7457), .Z(n7293) );
  AND U7356 ( .A(n10731), .B(n3593), .Z(n7457) );
  XOR U7357 ( .A(n7555), .B(n7556), .Z(n7290) );
  ANDN U7358 ( .A(n7557), .B(n7558), .Z(n7556) );
  XNOR U7359 ( .A(n7555), .B(n7559), .Z(n7557) );
  XOR U7360 ( .A(n7300), .B(n7560), .Z(n7294) );
  IV U7361 ( .A(n7299), .Z(n7560) );
  XNOR U7362 ( .A(n7296), .B(n7450), .Z(n7299) );
  AND U7363 ( .A(n11049), .B(n3166), .Z(n7450) );
  XOR U7364 ( .A(n7561), .B(n7562), .Z(n7296) );
  ANDN U7365 ( .A(n7563), .B(n7564), .Z(n7562) );
  XNOR U7366 ( .A(n7561), .B(n7565), .Z(n7563) );
  XOR U7367 ( .A(n7306), .B(n7566), .Z(n7300) );
  IV U7368 ( .A(n7305), .Z(n7566) );
  XNOR U7369 ( .A(n7302), .B(n7443), .Z(n7305) );
  AND U7370 ( .A(n11341), .B(n2765), .Z(n7443) );
  XOR U7371 ( .A(n7567), .B(n7568), .Z(n7302) );
  ANDN U7372 ( .A(n7569), .B(n7570), .Z(n7568) );
  XNOR U7373 ( .A(n7567), .B(n7571), .Z(n7569) );
  XOR U7374 ( .A(n7312), .B(n7572), .Z(n7306) );
  IV U7375 ( .A(n7311), .Z(n7572) );
  XNOR U7376 ( .A(n7308), .B(n7436), .Z(n7311) );
  AND U7377 ( .A(n11607), .B(n2396), .Z(n7436) );
  XOR U7378 ( .A(n7573), .B(n7574), .Z(n7308) );
  ANDN U7379 ( .A(n7575), .B(n7576), .Z(n7574) );
  XNOR U7380 ( .A(n7573), .B(n7577), .Z(n7575) );
  XOR U7381 ( .A(n7318), .B(n7578), .Z(n7312) );
  IV U7382 ( .A(n7317), .Z(n7578) );
  XNOR U7383 ( .A(n7314), .B(n7429), .Z(n7317) );
  AND U7384 ( .A(n11869), .B(n2053), .Z(n7429) );
  XOR U7385 ( .A(n7579), .B(n7580), .Z(n7314) );
  ANDN U7386 ( .A(n7581), .B(n7582), .Z(n7580) );
  XNOR U7387 ( .A(n7579), .B(n7583), .Z(n7581) );
  XOR U7388 ( .A(n7324), .B(n7584), .Z(n7318) );
  IV U7389 ( .A(n7323), .Z(n7584) );
  XNOR U7390 ( .A(n7320), .B(n7422), .Z(n7323) );
  AND U7391 ( .A(n12128), .B(n1737), .Z(n7422) );
  XOR U7392 ( .A(n7585), .B(n7586), .Z(n7320) );
  ANDN U7393 ( .A(n7587), .B(n7588), .Z(n7586) );
  XNOR U7394 ( .A(n7585), .B(n7589), .Z(n7587) );
  XOR U7395 ( .A(n7330), .B(n7590), .Z(n7324) );
  IV U7396 ( .A(n7329), .Z(n7590) );
  XNOR U7397 ( .A(n7326), .B(n7415), .Z(n7329) );
  AND U7398 ( .A(n12387), .B(n1448), .Z(n7415) );
  XOR U7399 ( .A(n7591), .B(n7592), .Z(n7326) );
  ANDN U7400 ( .A(n7593), .B(n7594), .Z(n7592) );
  XNOR U7401 ( .A(n7591), .B(n7595), .Z(n7593) );
  XOR U7402 ( .A(n7336), .B(n7596), .Z(n7330) );
  IV U7403 ( .A(n7335), .Z(n7596) );
  XNOR U7404 ( .A(n7332), .B(n7408), .Z(n7335) );
  AND U7405 ( .A(n12644), .B(n1185), .Z(n7408) );
  XOR U7406 ( .A(n7597), .B(n7598), .Z(n7332) );
  ANDN U7407 ( .A(n7599), .B(n7600), .Z(n7598) );
  XNOR U7408 ( .A(n7597), .B(n7601), .Z(n7599) );
  XOR U7409 ( .A(n7342), .B(n7602), .Z(n7336) );
  IV U7410 ( .A(n7341), .Z(n7602) );
  XNOR U7411 ( .A(n7338), .B(n7401), .Z(n7341) );
  AND U7412 ( .A(n12880), .B(n948), .Z(n7401) );
  XOR U7413 ( .A(n7603), .B(n7604), .Z(n7338) );
  ANDN U7414 ( .A(n7605), .B(n7606), .Z(n7604) );
  XNOR U7415 ( .A(n7603), .B(n7607), .Z(n7605) );
  XOR U7416 ( .A(n7348), .B(n7608), .Z(n7342) );
  IV U7417 ( .A(n7347), .Z(n7608) );
  XNOR U7418 ( .A(n7344), .B(n7394), .Z(n7347) );
  AND U7419 ( .A(n13070), .B(n736), .Z(n7394) );
  XOR U7420 ( .A(n7609), .B(n7610), .Z(n7344) );
  ANDN U7421 ( .A(n7611), .B(n7612), .Z(n7610) );
  XNOR U7422 ( .A(n7609), .B(n7613), .Z(n7611) );
  XOR U7423 ( .A(n7354), .B(n7614), .Z(n7348) );
  IV U7424 ( .A(n7353), .Z(n7614) );
  XNOR U7425 ( .A(n7350), .B(n7387), .Z(n7353) );
  AND U7426 ( .A(n13207), .B(n552), .Z(n7387) );
  XOR U7427 ( .A(n7615), .B(n7616), .Z(n7350) );
  ANDN U7428 ( .A(n7617), .B(n7618), .Z(n7616) );
  XNOR U7429 ( .A(n7615), .B(n7619), .Z(n7617) );
  XNOR U7430 ( .A(n7359), .B(n7112), .Z(n7354) );
  XNOR U7431 ( .A(n7356), .B(n7620), .Z(n7359) );
  AND U7432 ( .A(n6527), .B(n395), .Z(n7620) );
  XOR U7433 ( .A(n7621), .B(n7622), .Z(n7356) );
  ANDN U7434 ( .A(n7623), .B(n7624), .Z(n7622) );
  XNOR U7435 ( .A(n7384), .B(n7621), .Z(n7623) );
  XOR U7436 ( .A(n7625), .B(n7112), .Z(n7381) );
  NANDN U7437 ( .B(n6808), .A(n264), .Z(n7112) );
  XOR U7438 ( .A(n7626), .B(n7627), .Z(n264) );
  AND U7439 ( .A(n6809), .B(n7628), .Z(n7627) );
  XNOR U7440 ( .A(n7626), .B(n7366), .Z(n7628) );
  XOR U7441 ( .A(n7364), .B(n7626), .Z(n7366) );
  XOR U7442 ( .A(n7629), .B(n7630), .Z(n7364) );
  ANDN U7443 ( .A(n7629), .B(n7631), .Z(n7630) );
  XOR U7444 ( .A(n7632), .B(n7368), .Z(n7626) );
  IV U7445 ( .A(n7369), .Z(n7625) );
  XOR U7446 ( .A(n7633), .B(n7634), .Z(n7369) );
  AND U7447 ( .A(n7635), .B(n7636), .Z(n7634) );
  XOR U7448 ( .A(n7637), .B(n7633), .Z(n7636) );
  XOR U7449 ( .A(n7373), .B(n7377), .Z(n7380) );
  XOR U7450 ( .A(n7638), .B(n7639), .Z(n7373) );
  IV U7451 ( .A(n7640), .Z(n7639) );
  XOR U7452 ( .A(n7641), .B(n7642), .Z(n7377) );
  AND U7453 ( .A(n7641), .B(n7643), .Z(n7642) );
  XOR U7454 ( .A(n7644), .B(n7635), .Z(n7643) );
  XOR U7455 ( .A(n7645), .B(n7385), .Z(n7635) );
  XOR U7456 ( .A(n7392), .B(n7646), .Z(n7385) );
  IV U7457 ( .A(n7390), .Z(n7646) );
  XNOR U7458 ( .A(n7647), .B(n7389), .Z(n7390) );
  OR U7459 ( .A(n7648), .B(n7649), .Z(n7389) );
  NANDN U7460 ( .B(n6541), .A(n552), .Z(n7647) );
  XOR U7461 ( .A(n7399), .B(n7650), .Z(n7392) );
  IV U7462 ( .A(n7398), .Z(n7650) );
  XNOR U7463 ( .A(n7395), .B(n7651), .Z(n7398) );
  XOR U7464 ( .A(n7652), .B(n7653), .Z(n7395) );
  NANDN U7465 ( .B(n7654), .A(n7655), .Z(n7652) );
  XOR U7466 ( .A(n7653), .B(n7656), .Z(n7655) );
  XOR U7467 ( .A(n7406), .B(n7657), .Z(n7399) );
  IV U7468 ( .A(n7405), .Z(n7657) );
  XNOR U7469 ( .A(n7402), .B(n7658), .Z(n7405) );
  XOR U7470 ( .A(n7659), .B(n7660), .Z(n7402) );
  ANDN U7471 ( .A(n7661), .B(n7662), .Z(n7660) );
  XNOR U7472 ( .A(n7659), .B(n7663), .Z(n7661) );
  XOR U7473 ( .A(n7413), .B(n7664), .Z(n7406) );
  IV U7474 ( .A(n7412), .Z(n7664) );
  XNOR U7475 ( .A(n7409), .B(n7665), .Z(n7412) );
  XOR U7476 ( .A(n7666), .B(n7667), .Z(n7409) );
  ANDN U7477 ( .A(n7668), .B(n7669), .Z(n7667) );
  XNOR U7478 ( .A(n7666), .B(n7670), .Z(n7668) );
  XOR U7479 ( .A(n7420), .B(n7671), .Z(n7413) );
  IV U7480 ( .A(n7419), .Z(n7671) );
  XNOR U7481 ( .A(n7416), .B(n7672), .Z(n7419) );
  XOR U7482 ( .A(n7673), .B(n7674), .Z(n7416) );
  ANDN U7483 ( .A(n7675), .B(n7676), .Z(n7674) );
  XNOR U7484 ( .A(n7673), .B(n7677), .Z(n7675) );
  XOR U7485 ( .A(n7427), .B(n7678), .Z(n7420) );
  IV U7486 ( .A(n7426), .Z(n7678) );
  XNOR U7487 ( .A(n7423), .B(n7679), .Z(n7426) );
  XOR U7488 ( .A(n7680), .B(n7681), .Z(n7423) );
  ANDN U7489 ( .A(n7682), .B(n7683), .Z(n7681) );
  XNOR U7490 ( .A(n7680), .B(n7684), .Z(n7682) );
  XOR U7491 ( .A(n7434), .B(n7685), .Z(n7427) );
  IV U7492 ( .A(n7433), .Z(n7685) );
  XNOR U7493 ( .A(n7430), .B(n7686), .Z(n7433) );
  XOR U7494 ( .A(n7687), .B(n7688), .Z(n7430) );
  ANDN U7495 ( .A(n7689), .B(n7690), .Z(n7688) );
  XNOR U7496 ( .A(n7687), .B(n7691), .Z(n7689) );
  XOR U7497 ( .A(n7441), .B(n7692), .Z(n7434) );
  IV U7498 ( .A(n7440), .Z(n7692) );
  XNOR U7499 ( .A(n7437), .B(n7693), .Z(n7440) );
  XOR U7500 ( .A(n7694), .B(n7695), .Z(n7437) );
  ANDN U7501 ( .A(n7696), .B(n7697), .Z(n7695) );
  XNOR U7502 ( .A(n7694), .B(n7698), .Z(n7696) );
  XOR U7503 ( .A(n7448), .B(n7699), .Z(n7441) );
  IV U7504 ( .A(n7447), .Z(n7699) );
  XNOR U7505 ( .A(n7444), .B(n7700), .Z(n7447) );
  XOR U7506 ( .A(n7701), .B(n7702), .Z(n7444) );
  ANDN U7507 ( .A(n7703), .B(n7704), .Z(n7702) );
  XNOR U7508 ( .A(n7701), .B(n7705), .Z(n7703) );
  XOR U7509 ( .A(n7455), .B(n7706), .Z(n7448) );
  IV U7510 ( .A(n7454), .Z(n7706) );
  XNOR U7511 ( .A(n7451), .B(n7707), .Z(n7454) );
  XOR U7512 ( .A(n7708), .B(n7709), .Z(n7451) );
  ANDN U7513 ( .A(n7710), .B(n7711), .Z(n7709) );
  XNOR U7514 ( .A(n7708), .B(n7712), .Z(n7710) );
  XOR U7515 ( .A(n7462), .B(n7713), .Z(n7455) );
  IV U7516 ( .A(n7461), .Z(n7713) );
  XNOR U7517 ( .A(n7458), .B(n7714), .Z(n7461) );
  XOR U7518 ( .A(n7715), .B(n7716), .Z(n7458) );
  ANDN U7519 ( .A(n7717), .B(n7718), .Z(n7716) );
  XNOR U7520 ( .A(n7715), .B(n7719), .Z(n7717) );
  XOR U7521 ( .A(n7469), .B(n7720), .Z(n7462) );
  IV U7522 ( .A(n7468), .Z(n7720) );
  XNOR U7523 ( .A(n7465), .B(n7721), .Z(n7468) );
  XOR U7524 ( .A(n7722), .B(n7723), .Z(n7465) );
  ANDN U7525 ( .A(n7724), .B(n7725), .Z(n7723) );
  XNOR U7526 ( .A(n7722), .B(n7726), .Z(n7724) );
  XOR U7527 ( .A(n7476), .B(n7727), .Z(n7469) );
  IV U7528 ( .A(n7475), .Z(n7727) );
  XNOR U7529 ( .A(n7472), .B(n7728), .Z(n7475) );
  XOR U7530 ( .A(n7729), .B(n7730), .Z(n7472) );
  ANDN U7531 ( .A(n7731), .B(n7732), .Z(n7730) );
  XNOR U7532 ( .A(n7729), .B(n7733), .Z(n7731) );
  XOR U7533 ( .A(n7483), .B(n7734), .Z(n7476) );
  IV U7534 ( .A(n7482), .Z(n7734) );
  XNOR U7535 ( .A(n7479), .B(n7735), .Z(n7482) );
  XOR U7536 ( .A(n7736), .B(n7737), .Z(n7479) );
  ANDN U7537 ( .A(n7738), .B(n7739), .Z(n7737) );
  XNOR U7538 ( .A(n7736), .B(n7740), .Z(n7738) );
  XOR U7539 ( .A(n7490), .B(n7741), .Z(n7483) );
  IV U7540 ( .A(n7489), .Z(n7741) );
  XNOR U7541 ( .A(n7486), .B(n7742), .Z(n7489) );
  XOR U7542 ( .A(n7743), .B(n7744), .Z(n7486) );
  ANDN U7543 ( .A(n7745), .B(n7746), .Z(n7744) );
  XNOR U7544 ( .A(n7743), .B(n7747), .Z(n7745) );
  XOR U7545 ( .A(n7497), .B(n7748), .Z(n7490) );
  IV U7546 ( .A(n7496), .Z(n7748) );
  XNOR U7547 ( .A(n7493), .B(n7749), .Z(n7496) );
  XOR U7548 ( .A(n7750), .B(n7751), .Z(n7493) );
  ANDN U7549 ( .A(n7752), .B(n7753), .Z(n7751) );
  XNOR U7550 ( .A(n7750), .B(n7754), .Z(n7752) );
  XOR U7551 ( .A(n7504), .B(n7755), .Z(n7497) );
  IV U7552 ( .A(n7503), .Z(n7755) );
  XNOR U7553 ( .A(n7500), .B(n7756), .Z(n7503) );
  XOR U7554 ( .A(n7757), .B(n7758), .Z(n7500) );
  ANDN U7555 ( .A(n7759), .B(n7760), .Z(n7758) );
  XNOR U7556 ( .A(n7757), .B(n7761), .Z(n7759) );
  XOR U7557 ( .A(n7511), .B(n7762), .Z(n7504) );
  IV U7558 ( .A(n7510), .Z(n7762) );
  XNOR U7559 ( .A(n7507), .B(n7763), .Z(n7510) );
  XOR U7560 ( .A(n7764), .B(n7765), .Z(n7507) );
  ANDN U7561 ( .A(n7766), .B(n7767), .Z(n7765) );
  XNOR U7562 ( .A(n7764), .B(n7768), .Z(n7766) );
  XOR U7563 ( .A(n7517), .B(n7769), .Z(n7511) );
  IV U7564 ( .A(n7516), .Z(n7769) );
  XNOR U7565 ( .A(n7513), .B(n7770), .Z(n7516) );
  XOR U7566 ( .A(n7771), .B(n7772), .Z(n7513) );
  ANDN U7567 ( .A(n7773), .B(n7774), .Z(n7772) );
  XNOR U7568 ( .A(n7771), .B(n7775), .Z(n7773) );
  XOR U7569 ( .A(n7523), .B(n7776), .Z(n7517) );
  IV U7570 ( .A(n7522), .Z(n7776) );
  XNOR U7571 ( .A(n7519), .B(n7763), .Z(n7522) );
  AND U7572 ( .A(n8272), .B(n7241), .Z(n7763) );
  XOR U7573 ( .A(n7777), .B(n7778), .Z(n7519) );
  ANDN U7574 ( .A(n7779), .B(n7780), .Z(n7778) );
  XNOR U7575 ( .A(n7777), .B(n7781), .Z(n7779) );
  XOR U7576 ( .A(n7529), .B(n7782), .Z(n7523) );
  IV U7577 ( .A(n7528), .Z(n7782) );
  XNOR U7578 ( .A(n7525), .B(n7756), .Z(n7528) );
  AND U7579 ( .A(n8748), .B(n6688), .Z(n7756) );
  XOR U7580 ( .A(n7783), .B(n7784), .Z(n7525) );
  ANDN U7581 ( .A(n7785), .B(n7786), .Z(n7784) );
  XNOR U7582 ( .A(n7783), .B(n7787), .Z(n7785) );
  XOR U7583 ( .A(n7535), .B(n7788), .Z(n7529) );
  IV U7584 ( .A(n7534), .Z(n7788) );
  XNOR U7585 ( .A(n7531), .B(n7749), .Z(n7534) );
  AND U7586 ( .A(n9198), .B(n6118), .Z(n7749) );
  XOR U7587 ( .A(n7789), .B(n7790), .Z(n7531) );
  ANDN U7588 ( .A(n7791), .B(n7792), .Z(n7790) );
  XNOR U7589 ( .A(n7789), .B(n7793), .Z(n7791) );
  XOR U7590 ( .A(n7541), .B(n7794), .Z(n7535) );
  IV U7591 ( .A(n7540), .Z(n7794) );
  XNOR U7592 ( .A(n7537), .B(n7742), .Z(n7540) );
  AND U7593 ( .A(n9621), .B(n5561), .Z(n7742) );
  XOR U7594 ( .A(n7795), .B(n7796), .Z(n7537) );
  ANDN U7595 ( .A(n7797), .B(n7798), .Z(n7796) );
  XNOR U7596 ( .A(n7795), .B(n7799), .Z(n7797) );
  XOR U7597 ( .A(n7547), .B(n7800), .Z(n7541) );
  IV U7598 ( .A(n7546), .Z(n7800) );
  XNOR U7599 ( .A(n7543), .B(n7735), .Z(n7546) );
  AND U7600 ( .A(n10017), .B(n5030), .Z(n7735) );
  XOR U7601 ( .A(n7801), .B(n7802), .Z(n7543) );
  ANDN U7602 ( .A(n7803), .B(n7804), .Z(n7802) );
  XNOR U7603 ( .A(n7801), .B(n7805), .Z(n7803) );
  XOR U7604 ( .A(n7553), .B(n7806), .Z(n7547) );
  IV U7605 ( .A(n7552), .Z(n7806) );
  XNOR U7606 ( .A(n7549), .B(n7728), .Z(n7552) );
  AND U7607 ( .A(n10387), .B(n4525), .Z(n7728) );
  XOR U7608 ( .A(n7807), .B(n7808), .Z(n7549) );
  ANDN U7609 ( .A(n7809), .B(n7810), .Z(n7808) );
  XNOR U7610 ( .A(n7807), .B(n7811), .Z(n7809) );
  XOR U7611 ( .A(n7559), .B(n7812), .Z(n7553) );
  IV U7612 ( .A(n7558), .Z(n7812) );
  XNOR U7613 ( .A(n7555), .B(n7721), .Z(n7558) );
  AND U7614 ( .A(n10731), .B(n4046), .Z(n7721) );
  XOR U7615 ( .A(n7813), .B(n7814), .Z(n7555) );
  ANDN U7616 ( .A(n7815), .B(n7816), .Z(n7814) );
  XNOR U7617 ( .A(n7813), .B(n7817), .Z(n7815) );
  XOR U7618 ( .A(n7565), .B(n7818), .Z(n7559) );
  IV U7619 ( .A(n7564), .Z(n7818) );
  XNOR U7620 ( .A(n7561), .B(n7714), .Z(n7564) );
  AND U7621 ( .A(n11049), .B(n3593), .Z(n7714) );
  XOR U7622 ( .A(n7819), .B(n7820), .Z(n7561) );
  ANDN U7623 ( .A(n7821), .B(n7822), .Z(n7820) );
  XNOR U7624 ( .A(n7819), .B(n7823), .Z(n7821) );
  XOR U7625 ( .A(n7571), .B(n7824), .Z(n7565) );
  IV U7626 ( .A(n7570), .Z(n7824) );
  XNOR U7627 ( .A(n7567), .B(n7707), .Z(n7570) );
  AND U7628 ( .A(n11341), .B(n3166), .Z(n7707) );
  XOR U7629 ( .A(n7825), .B(n7826), .Z(n7567) );
  ANDN U7630 ( .A(n7827), .B(n7828), .Z(n7826) );
  XNOR U7631 ( .A(n7825), .B(n7829), .Z(n7827) );
  XOR U7632 ( .A(n7577), .B(n7830), .Z(n7571) );
  IV U7633 ( .A(n7576), .Z(n7830) );
  XNOR U7634 ( .A(n7573), .B(n7700), .Z(n7576) );
  AND U7635 ( .A(n11607), .B(n2765), .Z(n7700) );
  XOR U7636 ( .A(n7831), .B(n7832), .Z(n7573) );
  ANDN U7637 ( .A(n7833), .B(n7834), .Z(n7832) );
  XNOR U7638 ( .A(n7831), .B(n7835), .Z(n7833) );
  XOR U7639 ( .A(n7583), .B(n7836), .Z(n7577) );
  IV U7640 ( .A(n7582), .Z(n7836) );
  XNOR U7641 ( .A(n7579), .B(n7693), .Z(n7582) );
  AND U7642 ( .A(n11869), .B(n2396), .Z(n7693) );
  XOR U7643 ( .A(n7837), .B(n7838), .Z(n7579) );
  ANDN U7644 ( .A(n7839), .B(n7840), .Z(n7838) );
  XNOR U7645 ( .A(n7837), .B(n7841), .Z(n7839) );
  XOR U7646 ( .A(n7589), .B(n7842), .Z(n7583) );
  IV U7647 ( .A(n7588), .Z(n7842) );
  XNOR U7648 ( .A(n7585), .B(n7686), .Z(n7588) );
  AND U7649 ( .A(n12128), .B(n2053), .Z(n7686) );
  XOR U7650 ( .A(n7843), .B(n7844), .Z(n7585) );
  ANDN U7651 ( .A(n7845), .B(n7846), .Z(n7844) );
  XNOR U7652 ( .A(n7843), .B(n7847), .Z(n7845) );
  XOR U7653 ( .A(n7595), .B(n7848), .Z(n7589) );
  IV U7654 ( .A(n7594), .Z(n7848) );
  XNOR U7655 ( .A(n7591), .B(n7679), .Z(n7594) );
  AND U7656 ( .A(n12387), .B(n1737), .Z(n7679) );
  XOR U7657 ( .A(n7849), .B(n7850), .Z(n7591) );
  ANDN U7658 ( .A(n7851), .B(n7852), .Z(n7850) );
  XNOR U7659 ( .A(n7849), .B(n7853), .Z(n7851) );
  XOR U7660 ( .A(n7601), .B(n7854), .Z(n7595) );
  IV U7661 ( .A(n7600), .Z(n7854) );
  XNOR U7662 ( .A(n7597), .B(n7672), .Z(n7600) );
  AND U7663 ( .A(n12644), .B(n1448), .Z(n7672) );
  XOR U7664 ( .A(n7855), .B(n7856), .Z(n7597) );
  ANDN U7665 ( .A(n7857), .B(n7858), .Z(n7856) );
  XNOR U7666 ( .A(n7855), .B(n7859), .Z(n7857) );
  XOR U7667 ( .A(n7607), .B(n7860), .Z(n7601) );
  IV U7668 ( .A(n7606), .Z(n7860) );
  XNOR U7669 ( .A(n7603), .B(n7665), .Z(n7606) );
  AND U7670 ( .A(n12880), .B(n1185), .Z(n7665) );
  XOR U7671 ( .A(n7861), .B(n7862), .Z(n7603) );
  ANDN U7672 ( .A(n7863), .B(n7864), .Z(n7862) );
  XNOR U7673 ( .A(n7861), .B(n7865), .Z(n7863) );
  XOR U7674 ( .A(n7613), .B(n7866), .Z(n7607) );
  IV U7675 ( .A(n7612), .Z(n7866) );
  XNOR U7676 ( .A(n7609), .B(n7658), .Z(n7612) );
  AND U7677 ( .A(n13070), .B(n948), .Z(n7658) );
  XOR U7678 ( .A(n7867), .B(n7868), .Z(n7609) );
  ANDN U7679 ( .A(n7869), .B(n7870), .Z(n7868) );
  XNOR U7680 ( .A(n7867), .B(n7871), .Z(n7869) );
  XOR U7681 ( .A(n7619), .B(n7872), .Z(n7613) );
  IV U7682 ( .A(n7618), .Z(n7872) );
  XNOR U7683 ( .A(n7615), .B(n7651), .Z(n7618) );
  AND U7684 ( .A(n13207), .B(n736), .Z(n7651) );
  XOR U7685 ( .A(n7873), .B(n7874), .Z(n7615) );
  ANDN U7686 ( .A(n7875), .B(n7876), .Z(n7874) );
  XNOR U7687 ( .A(n7873), .B(n7877), .Z(n7875) );
  XNOR U7688 ( .A(n7624), .B(n7384), .Z(n7619) );
  XNOR U7689 ( .A(n7621), .B(n7878), .Z(n7624) );
  AND U7690 ( .A(n6527), .B(n552), .Z(n7878) );
  XOR U7691 ( .A(n7879), .B(n7880), .Z(n7621) );
  ANDN U7692 ( .A(n7881), .B(n7882), .Z(n7880) );
  XNOR U7693 ( .A(n7648), .B(n7879), .Z(n7881) );
  XOR U7694 ( .A(n7883), .B(n7384), .Z(n7645) );
  NANDN U7695 ( .B(n6808), .A(n395), .Z(n7384) );
  XOR U7696 ( .A(n7884), .B(n7885), .Z(n395) );
  AND U7697 ( .A(n6809), .B(n7886), .Z(n7885) );
  XNOR U7698 ( .A(n7884), .B(n7631), .Z(n7886) );
  XOR U7699 ( .A(n7629), .B(n7884), .Z(n7631) );
  XOR U7700 ( .A(n7887), .B(n7888), .Z(n7629) );
  ANDN U7701 ( .A(n7887), .B(n7889), .Z(n7888) );
  XOR U7702 ( .A(n7890), .B(n7368), .Z(n7884) );
  IV U7703 ( .A(n7633), .Z(n7883) );
  XOR U7704 ( .A(n7891), .B(n7892), .Z(n7633) );
  AND U7705 ( .A(n7893), .B(n7894), .Z(n7892) );
  XOR U7706 ( .A(n7895), .B(n7891), .Z(n7894) );
  XOR U7707 ( .A(n7637), .B(n7641), .Z(n7644) );
  XOR U7708 ( .A(n7896), .B(n7897), .Z(n7637) );
  IV U7709 ( .A(n7898), .Z(n7897) );
  XOR U7710 ( .A(n7899), .B(n7900), .Z(n7641) );
  AND U7711 ( .A(n7899), .B(n7901), .Z(n7900) );
  XOR U7712 ( .A(n7902), .B(n7893), .Z(n7901) );
  XOR U7713 ( .A(n7903), .B(n7649), .Z(n7893) );
  XOR U7714 ( .A(n7656), .B(n7904), .Z(n7649) );
  IV U7715 ( .A(n7654), .Z(n7904) );
  XNOR U7716 ( .A(n7905), .B(n7653), .Z(n7654) );
  OR U7717 ( .A(n7906), .B(n7907), .Z(n7653) );
  NANDN U7718 ( .B(n6541), .A(n736), .Z(n7905) );
  XOR U7719 ( .A(n7663), .B(n7908), .Z(n7656) );
  IV U7720 ( .A(n7662), .Z(n7908) );
  XNOR U7721 ( .A(n7659), .B(n7909), .Z(n7662) );
  XOR U7722 ( .A(n7910), .B(n7911), .Z(n7659) );
  NANDN U7723 ( .B(n7912), .A(n7913), .Z(n7910) );
  XOR U7724 ( .A(n7911), .B(n7914), .Z(n7913) );
  XOR U7725 ( .A(n7670), .B(n7915), .Z(n7663) );
  IV U7726 ( .A(n7669), .Z(n7915) );
  XNOR U7727 ( .A(n7666), .B(n7916), .Z(n7669) );
  XOR U7728 ( .A(n7917), .B(n7918), .Z(n7666) );
  ANDN U7729 ( .A(n7919), .B(n7920), .Z(n7918) );
  XNOR U7730 ( .A(n7917), .B(n7921), .Z(n7919) );
  XOR U7731 ( .A(n7677), .B(n7922), .Z(n7670) );
  IV U7732 ( .A(n7676), .Z(n7922) );
  XNOR U7733 ( .A(n7673), .B(n7923), .Z(n7676) );
  XOR U7734 ( .A(n7924), .B(n7925), .Z(n7673) );
  ANDN U7735 ( .A(n7926), .B(n7927), .Z(n7925) );
  XNOR U7736 ( .A(n7924), .B(n7928), .Z(n7926) );
  XOR U7737 ( .A(n7684), .B(n7929), .Z(n7677) );
  IV U7738 ( .A(n7683), .Z(n7929) );
  XNOR U7739 ( .A(n7680), .B(n7930), .Z(n7683) );
  XOR U7740 ( .A(n7931), .B(n7932), .Z(n7680) );
  ANDN U7741 ( .A(n7933), .B(n7934), .Z(n7932) );
  XNOR U7742 ( .A(n7931), .B(n7935), .Z(n7933) );
  XOR U7743 ( .A(n7691), .B(n7936), .Z(n7684) );
  IV U7744 ( .A(n7690), .Z(n7936) );
  XNOR U7745 ( .A(n7687), .B(n7937), .Z(n7690) );
  XOR U7746 ( .A(n7938), .B(n7939), .Z(n7687) );
  ANDN U7747 ( .A(n7940), .B(n7941), .Z(n7939) );
  XNOR U7748 ( .A(n7938), .B(n7942), .Z(n7940) );
  XOR U7749 ( .A(n7698), .B(n7943), .Z(n7691) );
  IV U7750 ( .A(n7697), .Z(n7943) );
  XNOR U7751 ( .A(n7694), .B(n7944), .Z(n7697) );
  XOR U7752 ( .A(n7945), .B(n7946), .Z(n7694) );
  ANDN U7753 ( .A(n7947), .B(n7948), .Z(n7946) );
  XNOR U7754 ( .A(n7945), .B(n7949), .Z(n7947) );
  XOR U7755 ( .A(n7705), .B(n7950), .Z(n7698) );
  IV U7756 ( .A(n7704), .Z(n7950) );
  XNOR U7757 ( .A(n7701), .B(n7951), .Z(n7704) );
  XOR U7758 ( .A(n7952), .B(n7953), .Z(n7701) );
  ANDN U7759 ( .A(n7954), .B(n7955), .Z(n7953) );
  XNOR U7760 ( .A(n7952), .B(n7956), .Z(n7954) );
  XOR U7761 ( .A(n7712), .B(n7957), .Z(n7705) );
  IV U7762 ( .A(n7711), .Z(n7957) );
  XNOR U7763 ( .A(n7708), .B(n7958), .Z(n7711) );
  XOR U7764 ( .A(n7959), .B(n7960), .Z(n7708) );
  ANDN U7765 ( .A(n7961), .B(n7962), .Z(n7960) );
  XNOR U7766 ( .A(n7959), .B(n7963), .Z(n7961) );
  XOR U7767 ( .A(n7719), .B(n7964), .Z(n7712) );
  IV U7768 ( .A(n7718), .Z(n7964) );
  XNOR U7769 ( .A(n7715), .B(n7965), .Z(n7718) );
  XOR U7770 ( .A(n7966), .B(n7967), .Z(n7715) );
  ANDN U7771 ( .A(n7968), .B(n7969), .Z(n7967) );
  XNOR U7772 ( .A(n7966), .B(n7970), .Z(n7968) );
  XOR U7773 ( .A(n7726), .B(n7971), .Z(n7719) );
  IV U7774 ( .A(n7725), .Z(n7971) );
  XNOR U7775 ( .A(n7722), .B(n7972), .Z(n7725) );
  XOR U7776 ( .A(n7973), .B(n7974), .Z(n7722) );
  ANDN U7777 ( .A(n7975), .B(n7976), .Z(n7974) );
  XNOR U7778 ( .A(n7973), .B(n7977), .Z(n7975) );
  XOR U7779 ( .A(n7733), .B(n7978), .Z(n7726) );
  IV U7780 ( .A(n7732), .Z(n7978) );
  XNOR U7781 ( .A(n7729), .B(n7979), .Z(n7732) );
  XOR U7782 ( .A(n7980), .B(n7981), .Z(n7729) );
  ANDN U7783 ( .A(n7982), .B(n7983), .Z(n7981) );
  XNOR U7784 ( .A(n7980), .B(n7984), .Z(n7982) );
  XOR U7785 ( .A(n7740), .B(n7985), .Z(n7733) );
  IV U7786 ( .A(n7739), .Z(n7985) );
  XNOR U7787 ( .A(n7736), .B(n7986), .Z(n7739) );
  XOR U7788 ( .A(n7987), .B(n7988), .Z(n7736) );
  ANDN U7789 ( .A(n7989), .B(n7990), .Z(n7988) );
  XNOR U7790 ( .A(n7987), .B(n7991), .Z(n7989) );
  XOR U7791 ( .A(n7747), .B(n7992), .Z(n7740) );
  IV U7792 ( .A(n7746), .Z(n7992) );
  XNOR U7793 ( .A(n7743), .B(n7993), .Z(n7746) );
  XOR U7794 ( .A(n7994), .B(n7995), .Z(n7743) );
  ANDN U7795 ( .A(n7996), .B(n7997), .Z(n7995) );
  XNOR U7796 ( .A(n7994), .B(n7998), .Z(n7996) );
  XOR U7797 ( .A(n7754), .B(n7999), .Z(n7747) );
  IV U7798 ( .A(n7753), .Z(n7999) );
  XNOR U7799 ( .A(n7750), .B(n8000), .Z(n7753) );
  XOR U7800 ( .A(n8001), .B(n8002), .Z(n7750) );
  ANDN U7801 ( .A(n8003), .B(n8004), .Z(n8002) );
  XNOR U7802 ( .A(n8001), .B(n8005), .Z(n8003) );
  XOR U7803 ( .A(n7761), .B(n8006), .Z(n7754) );
  IV U7804 ( .A(n7760), .Z(n8006) );
  XNOR U7805 ( .A(n7757), .B(n8007), .Z(n7760) );
  XOR U7806 ( .A(n8008), .B(n8009), .Z(n7757) );
  ANDN U7807 ( .A(n8010), .B(n8011), .Z(n8009) );
  XNOR U7808 ( .A(n8008), .B(n8012), .Z(n8010) );
  XOR U7809 ( .A(n7768), .B(n8013), .Z(n7761) );
  IV U7810 ( .A(n7767), .Z(n8013) );
  XNOR U7811 ( .A(n7764), .B(n8014), .Z(n7767) );
  XOR U7812 ( .A(n8015), .B(n8016), .Z(n7764) );
  ANDN U7813 ( .A(n8017), .B(n8018), .Z(n8016) );
  XNOR U7814 ( .A(n8015), .B(n8019), .Z(n8017) );
  XOR U7815 ( .A(n7775), .B(n8020), .Z(n7768) );
  IV U7816 ( .A(n7774), .Z(n8020) );
  XNOR U7817 ( .A(n7771), .B(n8021), .Z(n7774) );
  XOR U7818 ( .A(n8022), .B(n8023), .Z(n7771) );
  ANDN U7819 ( .A(n8024), .B(n8025), .Z(n8023) );
  XNOR U7820 ( .A(n8022), .B(n8026), .Z(n8024) );
  XOR U7821 ( .A(n7781), .B(n8027), .Z(n7775) );
  IV U7822 ( .A(n7780), .Z(n8027) );
  XNOR U7823 ( .A(n7777), .B(n8021), .Z(n7780) );
  AND U7824 ( .A(n8272), .B(n7770), .Z(n8021) );
  XOR U7825 ( .A(n8028), .B(n8029), .Z(n7777) );
  ANDN U7826 ( .A(n8030), .B(n8031), .Z(n8029) );
  XNOR U7827 ( .A(n8028), .B(n8032), .Z(n8030) );
  XOR U7828 ( .A(n7787), .B(n8033), .Z(n7781) );
  IV U7829 ( .A(n7786), .Z(n8033) );
  XNOR U7830 ( .A(n7783), .B(n8014), .Z(n7786) );
  AND U7831 ( .A(n8748), .B(n7241), .Z(n8014) );
  XOR U7832 ( .A(n8034), .B(n8035), .Z(n7783) );
  ANDN U7833 ( .A(n8036), .B(n8037), .Z(n8035) );
  XNOR U7834 ( .A(n8034), .B(n8038), .Z(n8036) );
  XOR U7835 ( .A(n7793), .B(n8039), .Z(n7787) );
  IV U7836 ( .A(n7792), .Z(n8039) );
  XNOR U7837 ( .A(n7789), .B(n8007), .Z(n7792) );
  AND U7838 ( .A(n9198), .B(n6688), .Z(n8007) );
  XOR U7839 ( .A(n8040), .B(n8041), .Z(n7789) );
  ANDN U7840 ( .A(n8042), .B(n8043), .Z(n8041) );
  XNOR U7841 ( .A(n8040), .B(n8044), .Z(n8042) );
  XOR U7842 ( .A(n7799), .B(n8045), .Z(n7793) );
  IV U7843 ( .A(n7798), .Z(n8045) );
  XNOR U7844 ( .A(n7795), .B(n8000), .Z(n7798) );
  AND U7845 ( .A(n9621), .B(n6118), .Z(n8000) );
  XOR U7846 ( .A(n8046), .B(n8047), .Z(n7795) );
  ANDN U7847 ( .A(n8048), .B(n8049), .Z(n8047) );
  XNOR U7848 ( .A(n8046), .B(n8050), .Z(n8048) );
  XOR U7849 ( .A(n7805), .B(n8051), .Z(n7799) );
  IV U7850 ( .A(n7804), .Z(n8051) );
  XNOR U7851 ( .A(n7801), .B(n7993), .Z(n7804) );
  AND U7852 ( .A(n10017), .B(n5561), .Z(n7993) );
  XOR U7853 ( .A(n8052), .B(n8053), .Z(n7801) );
  ANDN U7854 ( .A(n8054), .B(n8055), .Z(n8053) );
  XNOR U7855 ( .A(n8052), .B(n8056), .Z(n8054) );
  XOR U7856 ( .A(n7811), .B(n8057), .Z(n7805) );
  IV U7857 ( .A(n7810), .Z(n8057) );
  XNOR U7858 ( .A(n7807), .B(n7986), .Z(n7810) );
  AND U7859 ( .A(n10387), .B(n5030), .Z(n7986) );
  XOR U7860 ( .A(n8058), .B(n8059), .Z(n7807) );
  ANDN U7861 ( .A(n8060), .B(n8061), .Z(n8059) );
  XNOR U7862 ( .A(n8058), .B(n8062), .Z(n8060) );
  XOR U7863 ( .A(n7817), .B(n8063), .Z(n7811) );
  IV U7864 ( .A(n7816), .Z(n8063) );
  XNOR U7865 ( .A(n7813), .B(n7979), .Z(n7816) );
  AND U7866 ( .A(n10731), .B(n4525), .Z(n7979) );
  XOR U7867 ( .A(n8064), .B(n8065), .Z(n7813) );
  ANDN U7868 ( .A(n8066), .B(n8067), .Z(n8065) );
  XNOR U7869 ( .A(n8064), .B(n8068), .Z(n8066) );
  XOR U7870 ( .A(n7823), .B(n8069), .Z(n7817) );
  IV U7871 ( .A(n7822), .Z(n8069) );
  XNOR U7872 ( .A(n7819), .B(n7972), .Z(n7822) );
  AND U7873 ( .A(n11049), .B(n4046), .Z(n7972) );
  XOR U7874 ( .A(n8070), .B(n8071), .Z(n7819) );
  ANDN U7875 ( .A(n8072), .B(n8073), .Z(n8071) );
  XNOR U7876 ( .A(n8070), .B(n8074), .Z(n8072) );
  XOR U7877 ( .A(n7829), .B(n8075), .Z(n7823) );
  IV U7878 ( .A(n7828), .Z(n8075) );
  XNOR U7879 ( .A(n7825), .B(n7965), .Z(n7828) );
  AND U7880 ( .A(n11341), .B(n3593), .Z(n7965) );
  XOR U7881 ( .A(n8076), .B(n8077), .Z(n7825) );
  ANDN U7882 ( .A(n8078), .B(n8079), .Z(n8077) );
  XNOR U7883 ( .A(n8076), .B(n8080), .Z(n8078) );
  XOR U7884 ( .A(n7835), .B(n8081), .Z(n7829) );
  IV U7885 ( .A(n7834), .Z(n8081) );
  XNOR U7886 ( .A(n7831), .B(n7958), .Z(n7834) );
  AND U7887 ( .A(n11607), .B(n3166), .Z(n7958) );
  XOR U7888 ( .A(n8082), .B(n8083), .Z(n7831) );
  ANDN U7889 ( .A(n8084), .B(n8085), .Z(n8083) );
  XNOR U7890 ( .A(n8082), .B(n8086), .Z(n8084) );
  XOR U7891 ( .A(n7841), .B(n8087), .Z(n7835) );
  IV U7892 ( .A(n7840), .Z(n8087) );
  XNOR U7893 ( .A(n7837), .B(n7951), .Z(n7840) );
  AND U7894 ( .A(n11869), .B(n2765), .Z(n7951) );
  XOR U7895 ( .A(n8088), .B(n8089), .Z(n7837) );
  ANDN U7896 ( .A(n8090), .B(n8091), .Z(n8089) );
  XNOR U7897 ( .A(n8088), .B(n8092), .Z(n8090) );
  XOR U7898 ( .A(n7847), .B(n8093), .Z(n7841) );
  IV U7899 ( .A(n7846), .Z(n8093) );
  XNOR U7900 ( .A(n7843), .B(n7944), .Z(n7846) );
  AND U7901 ( .A(n12128), .B(n2396), .Z(n7944) );
  XOR U7902 ( .A(n8094), .B(n8095), .Z(n7843) );
  ANDN U7903 ( .A(n8096), .B(n8097), .Z(n8095) );
  XNOR U7904 ( .A(n8094), .B(n8098), .Z(n8096) );
  XOR U7905 ( .A(n7853), .B(n8099), .Z(n7847) );
  IV U7906 ( .A(n7852), .Z(n8099) );
  XNOR U7907 ( .A(n7849), .B(n7937), .Z(n7852) );
  AND U7908 ( .A(n12387), .B(n2053), .Z(n7937) );
  XOR U7909 ( .A(n8100), .B(n8101), .Z(n7849) );
  ANDN U7910 ( .A(n8102), .B(n8103), .Z(n8101) );
  XNOR U7911 ( .A(n8100), .B(n8104), .Z(n8102) );
  XOR U7912 ( .A(n7859), .B(n8105), .Z(n7853) );
  IV U7913 ( .A(n7858), .Z(n8105) );
  XNOR U7914 ( .A(n7855), .B(n7930), .Z(n7858) );
  AND U7915 ( .A(n12644), .B(n1737), .Z(n7930) );
  XOR U7916 ( .A(n8106), .B(n8107), .Z(n7855) );
  ANDN U7917 ( .A(n8108), .B(n8109), .Z(n8107) );
  XNOR U7918 ( .A(n8106), .B(n8110), .Z(n8108) );
  XOR U7919 ( .A(n7865), .B(n8111), .Z(n7859) );
  IV U7920 ( .A(n7864), .Z(n8111) );
  XNOR U7921 ( .A(n7861), .B(n7923), .Z(n7864) );
  AND U7922 ( .A(n12880), .B(n1448), .Z(n7923) );
  XOR U7923 ( .A(n8112), .B(n8113), .Z(n7861) );
  ANDN U7924 ( .A(n8114), .B(n8115), .Z(n8113) );
  XNOR U7925 ( .A(n8112), .B(n8116), .Z(n8114) );
  XOR U7926 ( .A(n7871), .B(n8117), .Z(n7865) );
  IV U7927 ( .A(n7870), .Z(n8117) );
  XNOR U7928 ( .A(n7867), .B(n7916), .Z(n7870) );
  AND U7929 ( .A(n13070), .B(n1185), .Z(n7916) );
  XOR U7930 ( .A(n8118), .B(n8119), .Z(n7867) );
  ANDN U7931 ( .A(n8120), .B(n8121), .Z(n8119) );
  XNOR U7932 ( .A(n8118), .B(n8122), .Z(n8120) );
  XOR U7933 ( .A(n7877), .B(n8123), .Z(n7871) );
  IV U7934 ( .A(n7876), .Z(n8123) );
  XNOR U7935 ( .A(n7873), .B(n7909), .Z(n7876) );
  AND U7936 ( .A(n13207), .B(n948), .Z(n7909) );
  XOR U7937 ( .A(n8124), .B(n8125), .Z(n7873) );
  ANDN U7938 ( .A(n8126), .B(n8127), .Z(n8125) );
  XNOR U7939 ( .A(n8124), .B(n8128), .Z(n8126) );
  XNOR U7940 ( .A(n7882), .B(n7648), .Z(n7877) );
  XNOR U7941 ( .A(n7879), .B(n8129), .Z(n7882) );
  AND U7942 ( .A(n6527), .B(n736), .Z(n8129) );
  XOR U7943 ( .A(n8130), .B(n8131), .Z(n7879) );
  ANDN U7944 ( .A(n8132), .B(n8133), .Z(n8131) );
  XNOR U7945 ( .A(n7906), .B(n8130), .Z(n8132) );
  XOR U7946 ( .A(n8134), .B(n7648), .Z(n7903) );
  NANDN U7947 ( .B(n6808), .A(n552), .Z(n7648) );
  XOR U7948 ( .A(n8135), .B(n8136), .Z(n552) );
  AND U7949 ( .A(n6809), .B(n8137), .Z(n8136) );
  XNOR U7950 ( .A(n8135), .B(n7889), .Z(n8137) );
  XOR U7951 ( .A(n7887), .B(n8135), .Z(n7889) );
  XOR U7952 ( .A(n8138), .B(n8139), .Z(n7887) );
  ANDN U7953 ( .A(n8138), .B(n8140), .Z(n8139) );
  XOR U7954 ( .A(n8141), .B(n7368), .Z(n8135) );
  IV U7955 ( .A(n7891), .Z(n8134) );
  XOR U7956 ( .A(n8142), .B(n8143), .Z(n7891) );
  AND U7957 ( .A(n8144), .B(n8145), .Z(n8143) );
  XOR U7958 ( .A(n8146), .B(n8142), .Z(n8145) );
  XOR U7959 ( .A(n7895), .B(n7899), .Z(n7902) );
  XOR U7960 ( .A(n8147), .B(n8148), .Z(n7895) );
  IV U7961 ( .A(n8149), .Z(n8148) );
  XOR U7962 ( .A(n8150), .B(n8151), .Z(n7899) );
  AND U7963 ( .A(n8150), .B(n8152), .Z(n8151) );
  XOR U7964 ( .A(n8153), .B(n8144), .Z(n8152) );
  XOR U7965 ( .A(n8154), .B(n7907), .Z(n8144) );
  XOR U7966 ( .A(n7914), .B(n8155), .Z(n7907) );
  IV U7967 ( .A(n7912), .Z(n8155) );
  XNOR U7968 ( .A(n8156), .B(n7911), .Z(n7912) );
  OR U7969 ( .A(n8157), .B(n8158), .Z(n7911) );
  NANDN U7970 ( .B(n6541), .A(n948), .Z(n8156) );
  XOR U7971 ( .A(n7921), .B(n8159), .Z(n7914) );
  IV U7972 ( .A(n7920), .Z(n8159) );
  XNOR U7973 ( .A(n7917), .B(n8160), .Z(n7920) );
  XOR U7974 ( .A(n8161), .B(n8162), .Z(n7917) );
  NANDN U7975 ( .B(n8163), .A(n8164), .Z(n8161) );
  XOR U7976 ( .A(n8162), .B(n8165), .Z(n8164) );
  XOR U7977 ( .A(n7928), .B(n8166), .Z(n7921) );
  IV U7978 ( .A(n7927), .Z(n8166) );
  XNOR U7979 ( .A(n7924), .B(n8167), .Z(n7927) );
  XOR U7980 ( .A(n8168), .B(n8169), .Z(n7924) );
  ANDN U7981 ( .A(n8170), .B(n8171), .Z(n8169) );
  XNOR U7982 ( .A(n8168), .B(n8172), .Z(n8170) );
  XOR U7983 ( .A(n7935), .B(n8173), .Z(n7928) );
  IV U7984 ( .A(n7934), .Z(n8173) );
  XNOR U7985 ( .A(n7931), .B(n8174), .Z(n7934) );
  XOR U7986 ( .A(n8175), .B(n8176), .Z(n7931) );
  ANDN U7987 ( .A(n8177), .B(n8178), .Z(n8176) );
  XNOR U7988 ( .A(n8175), .B(n8179), .Z(n8177) );
  XOR U7989 ( .A(n7942), .B(n8180), .Z(n7935) );
  IV U7990 ( .A(n7941), .Z(n8180) );
  XNOR U7991 ( .A(n7938), .B(n8181), .Z(n7941) );
  XOR U7992 ( .A(n8182), .B(n8183), .Z(n7938) );
  ANDN U7993 ( .A(n8184), .B(n8185), .Z(n8183) );
  XNOR U7994 ( .A(n8182), .B(n8186), .Z(n8184) );
  XOR U7995 ( .A(n7949), .B(n8187), .Z(n7942) );
  IV U7996 ( .A(n7948), .Z(n8187) );
  XNOR U7997 ( .A(n7945), .B(n8188), .Z(n7948) );
  XOR U7998 ( .A(n8189), .B(n8190), .Z(n7945) );
  ANDN U7999 ( .A(n8191), .B(n8192), .Z(n8190) );
  XNOR U8000 ( .A(n8189), .B(n8193), .Z(n8191) );
  XOR U8001 ( .A(n7956), .B(n8194), .Z(n7949) );
  IV U8002 ( .A(n7955), .Z(n8194) );
  XNOR U8003 ( .A(n7952), .B(n8195), .Z(n7955) );
  XOR U8004 ( .A(n8196), .B(n8197), .Z(n7952) );
  ANDN U8005 ( .A(n8198), .B(n8199), .Z(n8197) );
  XNOR U8006 ( .A(n8196), .B(n8200), .Z(n8198) );
  XOR U8007 ( .A(n7963), .B(n8201), .Z(n7956) );
  IV U8008 ( .A(n7962), .Z(n8201) );
  XNOR U8009 ( .A(n7959), .B(n8202), .Z(n7962) );
  XOR U8010 ( .A(n8203), .B(n8204), .Z(n7959) );
  ANDN U8011 ( .A(n8205), .B(n8206), .Z(n8204) );
  XNOR U8012 ( .A(n8203), .B(n8207), .Z(n8205) );
  XOR U8013 ( .A(n7970), .B(n8208), .Z(n7963) );
  IV U8014 ( .A(n7969), .Z(n8208) );
  XNOR U8015 ( .A(n7966), .B(n8209), .Z(n7969) );
  XOR U8016 ( .A(n8210), .B(n8211), .Z(n7966) );
  ANDN U8017 ( .A(n8212), .B(n8213), .Z(n8211) );
  XNOR U8018 ( .A(n8210), .B(n8214), .Z(n8212) );
  XOR U8019 ( .A(n7977), .B(n8215), .Z(n7970) );
  IV U8020 ( .A(n7976), .Z(n8215) );
  XNOR U8021 ( .A(n7973), .B(n8216), .Z(n7976) );
  XOR U8022 ( .A(n8217), .B(n8218), .Z(n7973) );
  ANDN U8023 ( .A(n8219), .B(n8220), .Z(n8218) );
  XNOR U8024 ( .A(n8217), .B(n8221), .Z(n8219) );
  XOR U8025 ( .A(n7984), .B(n8222), .Z(n7977) );
  IV U8026 ( .A(n7983), .Z(n8222) );
  XNOR U8027 ( .A(n7980), .B(n8223), .Z(n7983) );
  XOR U8028 ( .A(n8224), .B(n8225), .Z(n7980) );
  ANDN U8029 ( .A(n8226), .B(n8227), .Z(n8225) );
  XNOR U8030 ( .A(n8224), .B(n8228), .Z(n8226) );
  XOR U8031 ( .A(n7991), .B(n8229), .Z(n7984) );
  IV U8032 ( .A(n7990), .Z(n8229) );
  XNOR U8033 ( .A(n7987), .B(n8230), .Z(n7990) );
  XOR U8034 ( .A(n8231), .B(n8232), .Z(n7987) );
  ANDN U8035 ( .A(n8233), .B(n8234), .Z(n8232) );
  XNOR U8036 ( .A(n8231), .B(n8235), .Z(n8233) );
  XOR U8037 ( .A(n7998), .B(n8236), .Z(n7991) );
  IV U8038 ( .A(n7997), .Z(n8236) );
  XNOR U8039 ( .A(n7994), .B(n8237), .Z(n7997) );
  XOR U8040 ( .A(n8238), .B(n8239), .Z(n7994) );
  ANDN U8041 ( .A(n8240), .B(n8241), .Z(n8239) );
  XNOR U8042 ( .A(n8238), .B(n8242), .Z(n8240) );
  XOR U8043 ( .A(n8005), .B(n8243), .Z(n7998) );
  IV U8044 ( .A(n8004), .Z(n8243) );
  XNOR U8045 ( .A(n8001), .B(n8244), .Z(n8004) );
  XOR U8046 ( .A(n8245), .B(n8246), .Z(n8001) );
  ANDN U8047 ( .A(n8247), .B(n8248), .Z(n8246) );
  XNOR U8048 ( .A(n8245), .B(n8249), .Z(n8247) );
  XOR U8049 ( .A(n8012), .B(n8250), .Z(n8005) );
  IV U8050 ( .A(n8011), .Z(n8250) );
  XNOR U8051 ( .A(n8008), .B(n8251), .Z(n8011) );
  XOR U8052 ( .A(n8252), .B(n8253), .Z(n8008) );
  ANDN U8053 ( .A(n8254), .B(n8255), .Z(n8253) );
  XNOR U8054 ( .A(n8252), .B(n8256), .Z(n8254) );
  XOR U8055 ( .A(n8019), .B(n8257), .Z(n8012) );
  IV U8056 ( .A(n8018), .Z(n8257) );
  XNOR U8057 ( .A(n8015), .B(n8258), .Z(n8018) );
  XOR U8058 ( .A(n8259), .B(n8260), .Z(n8015) );
  ANDN U8059 ( .A(n8261), .B(n8262), .Z(n8260) );
  XNOR U8060 ( .A(n8259), .B(n8263), .Z(n8261) );
  XOR U8061 ( .A(n8026), .B(n8264), .Z(n8019) );
  IV U8062 ( .A(n8025), .Z(n8264) );
  XNOR U8063 ( .A(n8022), .B(n8265), .Z(n8025) );
  XOR U8064 ( .A(n8266), .B(n8267), .Z(n8022) );
  ANDN U8065 ( .A(n8268), .B(n8269), .Z(n8267) );
  XNOR U8066 ( .A(n8266), .B(n8270), .Z(n8268) );
  XOR U8067 ( .A(n8032), .B(n8271), .Z(n8026) );
  IV U8068 ( .A(n8031), .Z(n8271) );
  XNOR U8069 ( .A(n8028), .B(n8272), .Z(n8031) );
  XOR U8070 ( .A(n8273), .B(n8274), .Z(n8028) );
  ANDN U8071 ( .A(n8275), .B(n8276), .Z(n8274) );
  XNOR U8072 ( .A(n8273), .B(n8277), .Z(n8275) );
  XOR U8073 ( .A(n8038), .B(n8278), .Z(n8032) );
  IV U8074 ( .A(n8037), .Z(n8278) );
  XNOR U8075 ( .A(n8034), .B(n8265), .Z(n8037) );
  AND U8076 ( .A(n8748), .B(n7770), .Z(n8265) );
  XOR U8077 ( .A(n8279), .B(n8280), .Z(n8034) );
  ANDN U8078 ( .A(n8281), .B(n8282), .Z(n8280) );
  XNOR U8079 ( .A(n8279), .B(n8283), .Z(n8281) );
  XOR U8080 ( .A(n8044), .B(n8284), .Z(n8038) );
  IV U8081 ( .A(n8043), .Z(n8284) );
  XNOR U8082 ( .A(n8040), .B(n8258), .Z(n8043) );
  AND U8083 ( .A(n9198), .B(n7241), .Z(n8258) );
  XOR U8084 ( .A(n8285), .B(n8286), .Z(n8040) );
  ANDN U8085 ( .A(n8287), .B(n8288), .Z(n8286) );
  XNOR U8086 ( .A(n8285), .B(n8289), .Z(n8287) );
  XOR U8087 ( .A(n8050), .B(n8290), .Z(n8044) );
  IV U8088 ( .A(n8049), .Z(n8290) );
  XNOR U8089 ( .A(n8046), .B(n8251), .Z(n8049) );
  AND U8090 ( .A(n9621), .B(n6688), .Z(n8251) );
  XOR U8091 ( .A(n8291), .B(n8292), .Z(n8046) );
  ANDN U8092 ( .A(n8293), .B(n8294), .Z(n8292) );
  XNOR U8093 ( .A(n8291), .B(n8295), .Z(n8293) );
  XOR U8094 ( .A(n8056), .B(n8296), .Z(n8050) );
  IV U8095 ( .A(n8055), .Z(n8296) );
  XNOR U8096 ( .A(n8052), .B(n8244), .Z(n8055) );
  AND U8097 ( .A(n10017), .B(n6118), .Z(n8244) );
  XOR U8098 ( .A(n8297), .B(n8298), .Z(n8052) );
  ANDN U8099 ( .A(n8299), .B(n8300), .Z(n8298) );
  XNOR U8100 ( .A(n8297), .B(n8301), .Z(n8299) );
  XOR U8101 ( .A(n8062), .B(n8302), .Z(n8056) );
  IV U8102 ( .A(n8061), .Z(n8302) );
  XNOR U8103 ( .A(n8058), .B(n8237), .Z(n8061) );
  AND U8104 ( .A(n10387), .B(n5561), .Z(n8237) );
  XOR U8105 ( .A(n8303), .B(n8304), .Z(n8058) );
  ANDN U8106 ( .A(n8305), .B(n8306), .Z(n8304) );
  XNOR U8107 ( .A(n8303), .B(n8307), .Z(n8305) );
  XOR U8108 ( .A(n8068), .B(n8308), .Z(n8062) );
  IV U8109 ( .A(n8067), .Z(n8308) );
  XNOR U8110 ( .A(n8064), .B(n8230), .Z(n8067) );
  AND U8111 ( .A(n10731), .B(n5030), .Z(n8230) );
  XOR U8112 ( .A(n8309), .B(n8310), .Z(n8064) );
  ANDN U8113 ( .A(n8311), .B(n8312), .Z(n8310) );
  XNOR U8114 ( .A(n8309), .B(n8313), .Z(n8311) );
  XOR U8115 ( .A(n8074), .B(n8314), .Z(n8068) );
  IV U8116 ( .A(n8073), .Z(n8314) );
  XNOR U8117 ( .A(n8070), .B(n8223), .Z(n8073) );
  AND U8118 ( .A(n11049), .B(n4525), .Z(n8223) );
  XOR U8119 ( .A(n8315), .B(n8316), .Z(n8070) );
  ANDN U8120 ( .A(n8317), .B(n8318), .Z(n8316) );
  XNOR U8121 ( .A(n8315), .B(n8319), .Z(n8317) );
  XOR U8122 ( .A(n8080), .B(n8320), .Z(n8074) );
  IV U8123 ( .A(n8079), .Z(n8320) );
  XNOR U8124 ( .A(n8076), .B(n8216), .Z(n8079) );
  AND U8125 ( .A(n11341), .B(n4046), .Z(n8216) );
  XOR U8126 ( .A(n8321), .B(n8322), .Z(n8076) );
  ANDN U8127 ( .A(n8323), .B(n8324), .Z(n8322) );
  XNOR U8128 ( .A(n8321), .B(n8325), .Z(n8323) );
  XOR U8129 ( .A(n8086), .B(n8326), .Z(n8080) );
  IV U8130 ( .A(n8085), .Z(n8326) );
  XNOR U8131 ( .A(n8082), .B(n8209), .Z(n8085) );
  AND U8132 ( .A(n11607), .B(n3593), .Z(n8209) );
  XOR U8133 ( .A(n8327), .B(n8328), .Z(n8082) );
  ANDN U8134 ( .A(n8329), .B(n8330), .Z(n8328) );
  XNOR U8135 ( .A(n8327), .B(n8331), .Z(n8329) );
  XOR U8136 ( .A(n8092), .B(n8332), .Z(n8086) );
  IV U8137 ( .A(n8091), .Z(n8332) );
  XNOR U8138 ( .A(n8088), .B(n8202), .Z(n8091) );
  AND U8139 ( .A(n11869), .B(n3166), .Z(n8202) );
  XOR U8140 ( .A(n8333), .B(n8334), .Z(n8088) );
  ANDN U8141 ( .A(n8335), .B(n8336), .Z(n8334) );
  XNOR U8142 ( .A(n8333), .B(n8337), .Z(n8335) );
  XOR U8143 ( .A(n8098), .B(n8338), .Z(n8092) );
  IV U8144 ( .A(n8097), .Z(n8338) );
  XNOR U8145 ( .A(n8094), .B(n8195), .Z(n8097) );
  AND U8146 ( .A(n12128), .B(n2765), .Z(n8195) );
  XOR U8147 ( .A(n8339), .B(n8340), .Z(n8094) );
  ANDN U8148 ( .A(n8341), .B(n8342), .Z(n8340) );
  XNOR U8149 ( .A(n8339), .B(n8343), .Z(n8341) );
  XOR U8150 ( .A(n8104), .B(n8344), .Z(n8098) );
  IV U8151 ( .A(n8103), .Z(n8344) );
  XNOR U8152 ( .A(n8100), .B(n8188), .Z(n8103) );
  AND U8153 ( .A(n12387), .B(n2396), .Z(n8188) );
  XOR U8154 ( .A(n8345), .B(n8346), .Z(n8100) );
  ANDN U8155 ( .A(n8347), .B(n8348), .Z(n8346) );
  XNOR U8156 ( .A(n8345), .B(n8349), .Z(n8347) );
  XOR U8157 ( .A(n8110), .B(n8350), .Z(n8104) );
  IV U8158 ( .A(n8109), .Z(n8350) );
  XNOR U8159 ( .A(n8106), .B(n8181), .Z(n8109) );
  AND U8160 ( .A(n12644), .B(n2053), .Z(n8181) );
  XOR U8161 ( .A(n8351), .B(n8352), .Z(n8106) );
  ANDN U8162 ( .A(n8353), .B(n8354), .Z(n8352) );
  XNOR U8163 ( .A(n8351), .B(n8355), .Z(n8353) );
  XOR U8164 ( .A(n8116), .B(n8356), .Z(n8110) );
  IV U8165 ( .A(n8115), .Z(n8356) );
  XNOR U8166 ( .A(n8112), .B(n8174), .Z(n8115) );
  AND U8167 ( .A(n12880), .B(n1737), .Z(n8174) );
  XOR U8168 ( .A(n8357), .B(n8358), .Z(n8112) );
  ANDN U8169 ( .A(n8359), .B(n8360), .Z(n8358) );
  XNOR U8170 ( .A(n8357), .B(n8361), .Z(n8359) );
  XOR U8171 ( .A(n8122), .B(n8362), .Z(n8116) );
  IV U8172 ( .A(n8121), .Z(n8362) );
  XNOR U8173 ( .A(n8118), .B(n8167), .Z(n8121) );
  AND U8174 ( .A(n13070), .B(n1448), .Z(n8167) );
  XOR U8175 ( .A(n8363), .B(n8364), .Z(n8118) );
  ANDN U8176 ( .A(n8365), .B(n8366), .Z(n8364) );
  XNOR U8177 ( .A(n8363), .B(n8367), .Z(n8365) );
  XOR U8178 ( .A(n8128), .B(n8368), .Z(n8122) );
  IV U8179 ( .A(n8127), .Z(n8368) );
  XNOR U8180 ( .A(n8124), .B(n8160), .Z(n8127) );
  AND U8181 ( .A(n13207), .B(n1185), .Z(n8160) );
  XOR U8182 ( .A(n8369), .B(n8370), .Z(n8124) );
  ANDN U8183 ( .A(n8371), .B(n8372), .Z(n8370) );
  XNOR U8184 ( .A(n8369), .B(n8373), .Z(n8371) );
  XNOR U8185 ( .A(n8133), .B(n7906), .Z(n8128) );
  XNOR U8186 ( .A(n8130), .B(n8374), .Z(n8133) );
  AND U8187 ( .A(n6527), .B(n948), .Z(n8374) );
  XOR U8188 ( .A(n8375), .B(n8376), .Z(n8130) );
  ANDN U8189 ( .A(n8377), .B(n8378), .Z(n8376) );
  XNOR U8190 ( .A(n8157), .B(n8375), .Z(n8377) );
  XOR U8191 ( .A(n8379), .B(n7906), .Z(n8154) );
  NANDN U8192 ( .B(n6808), .A(n736), .Z(n7906) );
  XOR U8193 ( .A(n8380), .B(n8381), .Z(n736) );
  AND U8194 ( .A(n6809), .B(n8382), .Z(n8381) );
  XNOR U8195 ( .A(n8380), .B(n8140), .Z(n8382) );
  XOR U8196 ( .A(n8138), .B(n8380), .Z(n8140) );
  XOR U8197 ( .A(n8383), .B(n8384), .Z(n8138) );
  ANDN U8198 ( .A(n8383), .B(n8385), .Z(n8384) );
  XOR U8199 ( .A(n8386), .B(n7368), .Z(n8380) );
  IV U8200 ( .A(n8142), .Z(n8379) );
  XOR U8201 ( .A(n8387), .B(n8388), .Z(n8142) );
  AND U8202 ( .A(n8389), .B(n8390), .Z(n8388) );
  XOR U8203 ( .A(n8391), .B(n8387), .Z(n8390) );
  XOR U8204 ( .A(n8146), .B(n8150), .Z(n8153) );
  XOR U8205 ( .A(n8392), .B(n8393), .Z(n8146) );
  IV U8206 ( .A(n8394), .Z(n8393) );
  XOR U8207 ( .A(n8395), .B(n8396), .Z(n8150) );
  AND U8208 ( .A(n8395), .B(n8397), .Z(n8396) );
  XOR U8209 ( .A(n8398), .B(n8389), .Z(n8397) );
  XOR U8210 ( .A(n8399), .B(n8158), .Z(n8389) );
  XOR U8211 ( .A(n8165), .B(n8400), .Z(n8158) );
  IV U8212 ( .A(n8163), .Z(n8400) );
  XNOR U8213 ( .A(n8401), .B(n8162), .Z(n8163) );
  OR U8214 ( .A(n8402), .B(n8403), .Z(n8162) );
  NANDN U8215 ( .B(n6541), .A(n1185), .Z(n8401) );
  XOR U8216 ( .A(n8172), .B(n8404), .Z(n8165) );
  IV U8217 ( .A(n8171), .Z(n8404) );
  XNOR U8218 ( .A(n8168), .B(n8405), .Z(n8171) );
  XOR U8219 ( .A(n8406), .B(n8407), .Z(n8168) );
  NANDN U8220 ( .B(n8408), .A(n8409), .Z(n8406) );
  XOR U8221 ( .A(n8407), .B(n8410), .Z(n8409) );
  XOR U8222 ( .A(n8179), .B(n8411), .Z(n8172) );
  IV U8223 ( .A(n8178), .Z(n8411) );
  XNOR U8224 ( .A(n8175), .B(n8412), .Z(n8178) );
  XOR U8225 ( .A(n8413), .B(n8414), .Z(n8175) );
  ANDN U8226 ( .A(n8415), .B(n8416), .Z(n8414) );
  XNOR U8227 ( .A(n8413), .B(n8417), .Z(n8415) );
  XOR U8228 ( .A(n8186), .B(n8418), .Z(n8179) );
  IV U8229 ( .A(n8185), .Z(n8418) );
  XNOR U8230 ( .A(n8182), .B(n8419), .Z(n8185) );
  XOR U8231 ( .A(n8420), .B(n8421), .Z(n8182) );
  ANDN U8232 ( .A(n8422), .B(n8423), .Z(n8421) );
  XNOR U8233 ( .A(n8420), .B(n8424), .Z(n8422) );
  XOR U8234 ( .A(n8193), .B(n8425), .Z(n8186) );
  IV U8235 ( .A(n8192), .Z(n8425) );
  XNOR U8236 ( .A(n8189), .B(n8426), .Z(n8192) );
  XOR U8237 ( .A(n8427), .B(n8428), .Z(n8189) );
  ANDN U8238 ( .A(n8429), .B(n8430), .Z(n8428) );
  XNOR U8239 ( .A(n8427), .B(n8431), .Z(n8429) );
  XOR U8240 ( .A(n8200), .B(n8432), .Z(n8193) );
  IV U8241 ( .A(n8199), .Z(n8432) );
  XNOR U8242 ( .A(n8196), .B(n8433), .Z(n8199) );
  XOR U8243 ( .A(n8434), .B(n8435), .Z(n8196) );
  ANDN U8244 ( .A(n8436), .B(n8437), .Z(n8435) );
  XNOR U8245 ( .A(n8434), .B(n8438), .Z(n8436) );
  XOR U8246 ( .A(n8207), .B(n8439), .Z(n8200) );
  IV U8247 ( .A(n8206), .Z(n8439) );
  XNOR U8248 ( .A(n8203), .B(n8440), .Z(n8206) );
  XOR U8249 ( .A(n8441), .B(n8442), .Z(n8203) );
  ANDN U8250 ( .A(n8443), .B(n8444), .Z(n8442) );
  XNOR U8251 ( .A(n8441), .B(n8445), .Z(n8443) );
  XOR U8252 ( .A(n8214), .B(n8446), .Z(n8207) );
  IV U8253 ( .A(n8213), .Z(n8446) );
  XNOR U8254 ( .A(n8210), .B(n8447), .Z(n8213) );
  XOR U8255 ( .A(n8448), .B(n8449), .Z(n8210) );
  ANDN U8256 ( .A(n8450), .B(n8451), .Z(n8449) );
  XNOR U8257 ( .A(n8448), .B(n8452), .Z(n8450) );
  XOR U8258 ( .A(n8221), .B(n8453), .Z(n8214) );
  IV U8259 ( .A(n8220), .Z(n8453) );
  XNOR U8260 ( .A(n8217), .B(n8454), .Z(n8220) );
  XOR U8261 ( .A(n8455), .B(n8456), .Z(n8217) );
  ANDN U8262 ( .A(n8457), .B(n8458), .Z(n8456) );
  XNOR U8263 ( .A(n8455), .B(n8459), .Z(n8457) );
  XOR U8264 ( .A(n8228), .B(n8460), .Z(n8221) );
  IV U8265 ( .A(n8227), .Z(n8460) );
  XNOR U8266 ( .A(n8224), .B(n8461), .Z(n8227) );
  XOR U8267 ( .A(n8462), .B(n8463), .Z(n8224) );
  ANDN U8268 ( .A(n8464), .B(n8465), .Z(n8463) );
  XNOR U8269 ( .A(n8462), .B(n8466), .Z(n8464) );
  XOR U8270 ( .A(n8235), .B(n8467), .Z(n8228) );
  IV U8271 ( .A(n8234), .Z(n8467) );
  XNOR U8272 ( .A(n8231), .B(n8468), .Z(n8234) );
  XOR U8273 ( .A(n8469), .B(n8470), .Z(n8231) );
  ANDN U8274 ( .A(n8471), .B(n8472), .Z(n8470) );
  XNOR U8275 ( .A(n8469), .B(n8473), .Z(n8471) );
  XOR U8276 ( .A(n8242), .B(n8474), .Z(n8235) );
  IV U8277 ( .A(n8241), .Z(n8474) );
  XNOR U8278 ( .A(n8238), .B(n8475), .Z(n8241) );
  XOR U8279 ( .A(n8476), .B(n8477), .Z(n8238) );
  ANDN U8280 ( .A(n8478), .B(n8479), .Z(n8477) );
  XNOR U8281 ( .A(n8476), .B(n8480), .Z(n8478) );
  XOR U8282 ( .A(n8249), .B(n8481), .Z(n8242) );
  IV U8283 ( .A(n8248), .Z(n8481) );
  XNOR U8284 ( .A(n8245), .B(n8482), .Z(n8248) );
  XOR U8285 ( .A(n8483), .B(n8484), .Z(n8245) );
  ANDN U8286 ( .A(n8485), .B(n8486), .Z(n8484) );
  XNOR U8287 ( .A(n8483), .B(n8487), .Z(n8485) );
  XOR U8288 ( .A(n8256), .B(n8488), .Z(n8249) );
  IV U8289 ( .A(n8255), .Z(n8488) );
  XNOR U8290 ( .A(n8252), .B(n8489), .Z(n8255) );
  XOR U8291 ( .A(n8490), .B(n8491), .Z(n8252) );
  ANDN U8292 ( .A(n8492), .B(n8493), .Z(n8491) );
  XNOR U8293 ( .A(n8490), .B(n8494), .Z(n8492) );
  XOR U8294 ( .A(n8263), .B(n8495), .Z(n8256) );
  IV U8295 ( .A(n8262), .Z(n8495) );
  XNOR U8296 ( .A(n8259), .B(n8496), .Z(n8262) );
  XOR U8297 ( .A(n8497), .B(n8498), .Z(n8259) );
  ANDN U8298 ( .A(n8499), .B(n8500), .Z(n8498) );
  XNOR U8299 ( .A(n8497), .B(n8501), .Z(n8499) );
  XOR U8300 ( .A(n8270), .B(n8502), .Z(n8263) );
  IV U8301 ( .A(n8269), .Z(n8502) );
  XNOR U8302 ( .A(n8266), .B(n8503), .Z(n8269) );
  XOR U8303 ( .A(n8504), .B(n8505), .Z(n8266) );
  ANDN U8304 ( .A(n8506), .B(n8507), .Z(n8505) );
  XNOR U8305 ( .A(n8504), .B(n8508), .Z(n8506) );
  XOR U8306 ( .A(n8277), .B(n8509), .Z(n8270) );
  IV U8307 ( .A(n8276), .Z(n8509) );
  XNOR U8308 ( .A(n8273), .B(n8510), .Z(n8276) );
  XOR U8309 ( .A(n8511), .B(n8512), .Z(n8273) );
  ANDN U8310 ( .A(n8513), .B(n8514), .Z(n8512) );
  XNOR U8311 ( .A(n8511), .B(n8515), .Z(n8513) );
  XOR U8312 ( .A(n8283), .B(n8516), .Z(n8277) );
  IV U8313 ( .A(n8282), .Z(n8516) );
  XNOR U8314 ( .A(n8279), .B(n8510), .Z(n8282) );
  AND U8315 ( .A(n8748), .B(n8272), .Z(n8510) );
  XOR U8316 ( .A(n8517), .B(n8518), .Z(n8279) );
  ANDN U8317 ( .A(n8519), .B(n8520), .Z(n8518) );
  XNOR U8318 ( .A(n8517), .B(n8521), .Z(n8519) );
  XOR U8319 ( .A(n8289), .B(n8522), .Z(n8283) );
  IV U8320 ( .A(n8288), .Z(n8522) );
  XNOR U8321 ( .A(n8285), .B(n8503), .Z(n8288) );
  AND U8322 ( .A(n9198), .B(n7770), .Z(n8503) );
  XOR U8323 ( .A(n8523), .B(n8524), .Z(n8285) );
  ANDN U8324 ( .A(n8525), .B(n8526), .Z(n8524) );
  XNOR U8325 ( .A(n8523), .B(n8527), .Z(n8525) );
  XOR U8326 ( .A(n8295), .B(n8528), .Z(n8289) );
  IV U8327 ( .A(n8294), .Z(n8528) );
  XNOR U8328 ( .A(n8291), .B(n8496), .Z(n8294) );
  AND U8329 ( .A(n9621), .B(n7241), .Z(n8496) );
  XOR U8330 ( .A(n8529), .B(n8530), .Z(n8291) );
  ANDN U8331 ( .A(n8531), .B(n8532), .Z(n8530) );
  XNOR U8332 ( .A(n8529), .B(n8533), .Z(n8531) );
  XOR U8333 ( .A(n8301), .B(n8534), .Z(n8295) );
  IV U8334 ( .A(n8300), .Z(n8534) );
  XNOR U8335 ( .A(n8297), .B(n8489), .Z(n8300) );
  AND U8336 ( .A(n10017), .B(n6688), .Z(n8489) );
  XOR U8337 ( .A(n8535), .B(n8536), .Z(n8297) );
  ANDN U8338 ( .A(n8537), .B(n8538), .Z(n8536) );
  XNOR U8339 ( .A(n8535), .B(n8539), .Z(n8537) );
  XOR U8340 ( .A(n8307), .B(n8540), .Z(n8301) );
  IV U8341 ( .A(n8306), .Z(n8540) );
  XNOR U8342 ( .A(n8303), .B(n8482), .Z(n8306) );
  AND U8343 ( .A(n10387), .B(n6118), .Z(n8482) );
  XOR U8344 ( .A(n8541), .B(n8542), .Z(n8303) );
  ANDN U8345 ( .A(n8543), .B(n8544), .Z(n8542) );
  XNOR U8346 ( .A(n8541), .B(n8545), .Z(n8543) );
  XOR U8347 ( .A(n8313), .B(n8546), .Z(n8307) );
  IV U8348 ( .A(n8312), .Z(n8546) );
  XNOR U8349 ( .A(n8309), .B(n8475), .Z(n8312) );
  AND U8350 ( .A(n10731), .B(n5561), .Z(n8475) );
  XOR U8351 ( .A(n8547), .B(n8548), .Z(n8309) );
  ANDN U8352 ( .A(n8549), .B(n8550), .Z(n8548) );
  XNOR U8353 ( .A(n8547), .B(n8551), .Z(n8549) );
  XOR U8354 ( .A(n8319), .B(n8552), .Z(n8313) );
  IV U8355 ( .A(n8318), .Z(n8552) );
  XNOR U8356 ( .A(n8315), .B(n8468), .Z(n8318) );
  AND U8357 ( .A(n11049), .B(n5030), .Z(n8468) );
  XOR U8358 ( .A(n8553), .B(n8554), .Z(n8315) );
  ANDN U8359 ( .A(n8555), .B(n8556), .Z(n8554) );
  XNOR U8360 ( .A(n8553), .B(n8557), .Z(n8555) );
  XOR U8361 ( .A(n8325), .B(n8558), .Z(n8319) );
  IV U8362 ( .A(n8324), .Z(n8558) );
  XNOR U8363 ( .A(n8321), .B(n8461), .Z(n8324) );
  AND U8364 ( .A(n11341), .B(n4525), .Z(n8461) );
  XOR U8365 ( .A(n8559), .B(n8560), .Z(n8321) );
  ANDN U8366 ( .A(n8561), .B(n8562), .Z(n8560) );
  XNOR U8367 ( .A(n8559), .B(n8563), .Z(n8561) );
  XOR U8368 ( .A(n8331), .B(n8564), .Z(n8325) );
  IV U8369 ( .A(n8330), .Z(n8564) );
  XNOR U8370 ( .A(n8327), .B(n8454), .Z(n8330) );
  AND U8371 ( .A(n11607), .B(n4046), .Z(n8454) );
  XOR U8372 ( .A(n8565), .B(n8566), .Z(n8327) );
  ANDN U8373 ( .A(n8567), .B(n8568), .Z(n8566) );
  XNOR U8374 ( .A(n8565), .B(n8569), .Z(n8567) );
  XOR U8375 ( .A(n8337), .B(n8570), .Z(n8331) );
  IV U8376 ( .A(n8336), .Z(n8570) );
  XNOR U8377 ( .A(n8333), .B(n8447), .Z(n8336) );
  AND U8378 ( .A(n11869), .B(n3593), .Z(n8447) );
  XOR U8379 ( .A(n8571), .B(n8572), .Z(n8333) );
  ANDN U8380 ( .A(n8573), .B(n8574), .Z(n8572) );
  XNOR U8381 ( .A(n8571), .B(n8575), .Z(n8573) );
  XOR U8382 ( .A(n8343), .B(n8576), .Z(n8337) );
  IV U8383 ( .A(n8342), .Z(n8576) );
  XNOR U8384 ( .A(n8339), .B(n8440), .Z(n8342) );
  AND U8385 ( .A(n12128), .B(n3166), .Z(n8440) );
  XOR U8386 ( .A(n8577), .B(n8578), .Z(n8339) );
  ANDN U8387 ( .A(n8579), .B(n8580), .Z(n8578) );
  XNOR U8388 ( .A(n8577), .B(n8581), .Z(n8579) );
  XOR U8389 ( .A(n8349), .B(n8582), .Z(n8343) );
  IV U8390 ( .A(n8348), .Z(n8582) );
  XNOR U8391 ( .A(n8345), .B(n8433), .Z(n8348) );
  AND U8392 ( .A(n12387), .B(n2765), .Z(n8433) );
  XOR U8393 ( .A(n8583), .B(n8584), .Z(n8345) );
  ANDN U8394 ( .A(n8585), .B(n8586), .Z(n8584) );
  XNOR U8395 ( .A(n8583), .B(n8587), .Z(n8585) );
  XOR U8396 ( .A(n8355), .B(n8588), .Z(n8349) );
  IV U8397 ( .A(n8354), .Z(n8588) );
  XNOR U8398 ( .A(n8351), .B(n8426), .Z(n8354) );
  AND U8399 ( .A(n12644), .B(n2396), .Z(n8426) );
  XOR U8400 ( .A(n8589), .B(n8590), .Z(n8351) );
  ANDN U8401 ( .A(n8591), .B(n8592), .Z(n8590) );
  XNOR U8402 ( .A(n8589), .B(n8593), .Z(n8591) );
  XOR U8403 ( .A(n8361), .B(n8594), .Z(n8355) );
  IV U8404 ( .A(n8360), .Z(n8594) );
  XNOR U8405 ( .A(n8357), .B(n8419), .Z(n8360) );
  AND U8406 ( .A(n12880), .B(n2053), .Z(n8419) );
  XOR U8407 ( .A(n8595), .B(n8596), .Z(n8357) );
  ANDN U8408 ( .A(n8597), .B(n8598), .Z(n8596) );
  XNOR U8409 ( .A(n8595), .B(n8599), .Z(n8597) );
  XOR U8410 ( .A(n8367), .B(n8600), .Z(n8361) );
  IV U8411 ( .A(n8366), .Z(n8600) );
  XNOR U8412 ( .A(n8363), .B(n8412), .Z(n8366) );
  AND U8413 ( .A(n13070), .B(n1737), .Z(n8412) );
  XOR U8414 ( .A(n8601), .B(n8602), .Z(n8363) );
  ANDN U8415 ( .A(n8603), .B(n8604), .Z(n8602) );
  XNOR U8416 ( .A(n8601), .B(n8605), .Z(n8603) );
  XOR U8417 ( .A(n8373), .B(n8606), .Z(n8367) );
  IV U8418 ( .A(n8372), .Z(n8606) );
  XNOR U8419 ( .A(n8369), .B(n8405), .Z(n8372) );
  AND U8420 ( .A(n13207), .B(n1448), .Z(n8405) );
  XOR U8421 ( .A(n8607), .B(n8608), .Z(n8369) );
  ANDN U8422 ( .A(n8609), .B(n8610), .Z(n8608) );
  XNOR U8423 ( .A(n8607), .B(n8611), .Z(n8609) );
  XNOR U8424 ( .A(n8378), .B(n8157), .Z(n8373) );
  XNOR U8425 ( .A(n8375), .B(n8612), .Z(n8378) );
  AND U8426 ( .A(n6527), .B(n1185), .Z(n8612) );
  XOR U8427 ( .A(n8613), .B(n8614), .Z(n8375) );
  ANDN U8428 ( .A(n8615), .B(n8616), .Z(n8614) );
  XNOR U8429 ( .A(n8402), .B(n8613), .Z(n8615) );
  XOR U8430 ( .A(n8617), .B(n8157), .Z(n8399) );
  NANDN U8431 ( .B(n6808), .A(n948), .Z(n8157) );
  XOR U8432 ( .A(n8618), .B(n8619), .Z(n948) );
  AND U8433 ( .A(n6809), .B(n8620), .Z(n8619) );
  XNOR U8434 ( .A(n8618), .B(n8385), .Z(n8620) );
  XOR U8435 ( .A(n8383), .B(n8618), .Z(n8385) );
  XOR U8436 ( .A(n8621), .B(n8622), .Z(n8383) );
  ANDN U8437 ( .A(n8621), .B(n8623), .Z(n8622) );
  XOR U8438 ( .A(n8624), .B(n7368), .Z(n8618) );
  IV U8439 ( .A(n8387), .Z(n8617) );
  XOR U8440 ( .A(n8625), .B(n8626), .Z(n8387) );
  AND U8441 ( .A(n8627), .B(n8628), .Z(n8626) );
  XOR U8442 ( .A(n8629), .B(n8625), .Z(n8628) );
  XOR U8443 ( .A(n8391), .B(n8395), .Z(n8398) );
  XOR U8444 ( .A(n8630), .B(n8631), .Z(n8391) );
  IV U8445 ( .A(n8632), .Z(n8631) );
  XOR U8446 ( .A(n8633), .B(n8634), .Z(n8395) );
  AND U8447 ( .A(n8633), .B(n8635), .Z(n8634) );
  XOR U8448 ( .A(n8636), .B(n8627), .Z(n8635) );
  XOR U8449 ( .A(n8637), .B(n8403), .Z(n8627) );
  XOR U8450 ( .A(n8410), .B(n8638), .Z(n8403) );
  IV U8451 ( .A(n8408), .Z(n8638) );
  XNOR U8452 ( .A(n8639), .B(n8407), .Z(n8408) );
  OR U8453 ( .A(n8640), .B(n8641), .Z(n8407) );
  NANDN U8454 ( .B(n6541), .A(n1448), .Z(n8639) );
  XOR U8455 ( .A(n8417), .B(n8642), .Z(n8410) );
  IV U8456 ( .A(n8416), .Z(n8642) );
  XNOR U8457 ( .A(n8413), .B(n8643), .Z(n8416) );
  XOR U8458 ( .A(n8644), .B(n8645), .Z(n8413) );
  NANDN U8459 ( .B(n8646), .A(n8647), .Z(n8644) );
  XOR U8460 ( .A(n8645), .B(n8648), .Z(n8647) );
  XOR U8461 ( .A(n8424), .B(n8649), .Z(n8417) );
  IV U8462 ( .A(n8423), .Z(n8649) );
  XNOR U8463 ( .A(n8420), .B(n8650), .Z(n8423) );
  XOR U8464 ( .A(n8651), .B(n8652), .Z(n8420) );
  ANDN U8465 ( .A(n8653), .B(n8654), .Z(n8652) );
  XNOR U8466 ( .A(n8651), .B(n8655), .Z(n8653) );
  XOR U8467 ( .A(n8431), .B(n8656), .Z(n8424) );
  IV U8468 ( .A(n8430), .Z(n8656) );
  XNOR U8469 ( .A(n8427), .B(n8657), .Z(n8430) );
  XOR U8470 ( .A(n8658), .B(n8659), .Z(n8427) );
  ANDN U8471 ( .A(n8660), .B(n8661), .Z(n8659) );
  XNOR U8472 ( .A(n8658), .B(n8662), .Z(n8660) );
  XOR U8473 ( .A(n8438), .B(n8663), .Z(n8431) );
  IV U8474 ( .A(n8437), .Z(n8663) );
  XNOR U8475 ( .A(n8434), .B(n8664), .Z(n8437) );
  XOR U8476 ( .A(n8665), .B(n8666), .Z(n8434) );
  ANDN U8477 ( .A(n8667), .B(n8668), .Z(n8666) );
  XNOR U8478 ( .A(n8665), .B(n8669), .Z(n8667) );
  XOR U8479 ( .A(n8445), .B(n8670), .Z(n8438) );
  IV U8480 ( .A(n8444), .Z(n8670) );
  XNOR U8481 ( .A(n8441), .B(n8671), .Z(n8444) );
  XOR U8482 ( .A(n8672), .B(n8673), .Z(n8441) );
  ANDN U8483 ( .A(n8674), .B(n8675), .Z(n8673) );
  XNOR U8484 ( .A(n8672), .B(n8676), .Z(n8674) );
  XOR U8485 ( .A(n8452), .B(n8677), .Z(n8445) );
  IV U8486 ( .A(n8451), .Z(n8677) );
  XNOR U8487 ( .A(n8448), .B(n8678), .Z(n8451) );
  XOR U8488 ( .A(n8679), .B(n8680), .Z(n8448) );
  ANDN U8489 ( .A(n8681), .B(n8682), .Z(n8680) );
  XNOR U8490 ( .A(n8679), .B(n8683), .Z(n8681) );
  XOR U8491 ( .A(n8459), .B(n8684), .Z(n8452) );
  IV U8492 ( .A(n8458), .Z(n8684) );
  XNOR U8493 ( .A(n8455), .B(n8685), .Z(n8458) );
  XOR U8494 ( .A(n8686), .B(n8687), .Z(n8455) );
  ANDN U8495 ( .A(n8688), .B(n8689), .Z(n8687) );
  XNOR U8496 ( .A(n8686), .B(n8690), .Z(n8688) );
  XOR U8497 ( .A(n8466), .B(n8691), .Z(n8459) );
  IV U8498 ( .A(n8465), .Z(n8691) );
  XNOR U8499 ( .A(n8462), .B(n8692), .Z(n8465) );
  XOR U8500 ( .A(n8693), .B(n8694), .Z(n8462) );
  ANDN U8501 ( .A(n8695), .B(n8696), .Z(n8694) );
  XNOR U8502 ( .A(n8693), .B(n8697), .Z(n8695) );
  XOR U8503 ( .A(n8473), .B(n8698), .Z(n8466) );
  IV U8504 ( .A(n8472), .Z(n8698) );
  XNOR U8505 ( .A(n8469), .B(n8699), .Z(n8472) );
  XOR U8506 ( .A(n8700), .B(n8701), .Z(n8469) );
  ANDN U8507 ( .A(n8702), .B(n8703), .Z(n8701) );
  XNOR U8508 ( .A(n8700), .B(n8704), .Z(n8702) );
  XOR U8509 ( .A(n8480), .B(n8705), .Z(n8473) );
  IV U8510 ( .A(n8479), .Z(n8705) );
  XNOR U8511 ( .A(n8476), .B(n8706), .Z(n8479) );
  XOR U8512 ( .A(n8707), .B(n8708), .Z(n8476) );
  ANDN U8513 ( .A(n8709), .B(n8710), .Z(n8708) );
  XNOR U8514 ( .A(n8707), .B(n8711), .Z(n8709) );
  XOR U8515 ( .A(n8487), .B(n8712), .Z(n8480) );
  IV U8516 ( .A(n8486), .Z(n8712) );
  XNOR U8517 ( .A(n8483), .B(n8713), .Z(n8486) );
  XOR U8518 ( .A(n8714), .B(n8715), .Z(n8483) );
  ANDN U8519 ( .A(n8716), .B(n8717), .Z(n8715) );
  XNOR U8520 ( .A(n8714), .B(n8718), .Z(n8716) );
  XOR U8521 ( .A(n8494), .B(n8719), .Z(n8487) );
  IV U8522 ( .A(n8493), .Z(n8719) );
  XNOR U8523 ( .A(n8490), .B(n8720), .Z(n8493) );
  XOR U8524 ( .A(n8721), .B(n8722), .Z(n8490) );
  ANDN U8525 ( .A(n8723), .B(n8724), .Z(n8722) );
  XNOR U8526 ( .A(n8721), .B(n8725), .Z(n8723) );
  XOR U8527 ( .A(n8501), .B(n8726), .Z(n8494) );
  IV U8528 ( .A(n8500), .Z(n8726) );
  XNOR U8529 ( .A(n8497), .B(n8727), .Z(n8500) );
  XOR U8530 ( .A(n8728), .B(n8729), .Z(n8497) );
  ANDN U8531 ( .A(n8730), .B(n8731), .Z(n8729) );
  XNOR U8532 ( .A(n8728), .B(n8732), .Z(n8730) );
  XOR U8533 ( .A(n8508), .B(n8733), .Z(n8501) );
  IV U8534 ( .A(n8507), .Z(n8733) );
  XNOR U8535 ( .A(n8504), .B(n8734), .Z(n8507) );
  XOR U8536 ( .A(n8735), .B(n8736), .Z(n8504) );
  ANDN U8537 ( .A(n8737), .B(n8738), .Z(n8736) );
  XNOR U8538 ( .A(n8735), .B(n8739), .Z(n8737) );
  XOR U8539 ( .A(n8515), .B(n8740), .Z(n8508) );
  IV U8540 ( .A(n8514), .Z(n8740) );
  XNOR U8541 ( .A(n8511), .B(n8741), .Z(n8514) );
  XOR U8542 ( .A(n8742), .B(n8743), .Z(n8511) );
  ANDN U8543 ( .A(n8744), .B(n8745), .Z(n8743) );
  XNOR U8544 ( .A(n8742), .B(n8746), .Z(n8744) );
  XOR U8545 ( .A(n8521), .B(n8747), .Z(n8515) );
  IV U8546 ( .A(n8520), .Z(n8747) );
  XNOR U8547 ( .A(n8517), .B(n8748), .Z(n8520) );
  XOR U8548 ( .A(n8749), .B(n8750), .Z(n8517) );
  ANDN U8549 ( .A(n8751), .B(n8752), .Z(n8750) );
  XNOR U8550 ( .A(n8749), .B(n8753), .Z(n8751) );
  XOR U8551 ( .A(n8527), .B(n8754), .Z(n8521) );
  IV U8552 ( .A(n8526), .Z(n8754) );
  XNOR U8553 ( .A(n8523), .B(n8741), .Z(n8526) );
  AND U8554 ( .A(n9198), .B(n8272), .Z(n8741) );
  XOR U8555 ( .A(n8755), .B(n8756), .Z(n8523) );
  ANDN U8556 ( .A(n8757), .B(n8758), .Z(n8756) );
  XNOR U8557 ( .A(n8755), .B(n8759), .Z(n8757) );
  XOR U8558 ( .A(n8533), .B(n8760), .Z(n8527) );
  IV U8559 ( .A(n8532), .Z(n8760) );
  XNOR U8560 ( .A(n8529), .B(n8734), .Z(n8532) );
  AND U8561 ( .A(n9621), .B(n7770), .Z(n8734) );
  XOR U8562 ( .A(n8761), .B(n8762), .Z(n8529) );
  ANDN U8563 ( .A(n8763), .B(n8764), .Z(n8762) );
  XNOR U8564 ( .A(n8761), .B(n8765), .Z(n8763) );
  XOR U8565 ( .A(n8539), .B(n8766), .Z(n8533) );
  IV U8566 ( .A(n8538), .Z(n8766) );
  XNOR U8567 ( .A(n8535), .B(n8727), .Z(n8538) );
  AND U8568 ( .A(n10017), .B(n7241), .Z(n8727) );
  XOR U8569 ( .A(n8767), .B(n8768), .Z(n8535) );
  ANDN U8570 ( .A(n8769), .B(n8770), .Z(n8768) );
  XNOR U8571 ( .A(n8767), .B(n8771), .Z(n8769) );
  XOR U8572 ( .A(n8545), .B(n8772), .Z(n8539) );
  IV U8573 ( .A(n8544), .Z(n8772) );
  XNOR U8574 ( .A(n8541), .B(n8720), .Z(n8544) );
  AND U8575 ( .A(n10387), .B(n6688), .Z(n8720) );
  XOR U8576 ( .A(n8773), .B(n8774), .Z(n8541) );
  ANDN U8577 ( .A(n8775), .B(n8776), .Z(n8774) );
  XNOR U8578 ( .A(n8773), .B(n8777), .Z(n8775) );
  XOR U8579 ( .A(n8551), .B(n8778), .Z(n8545) );
  IV U8580 ( .A(n8550), .Z(n8778) );
  XNOR U8581 ( .A(n8547), .B(n8713), .Z(n8550) );
  AND U8582 ( .A(n10731), .B(n6118), .Z(n8713) );
  XOR U8583 ( .A(n8779), .B(n8780), .Z(n8547) );
  ANDN U8584 ( .A(n8781), .B(n8782), .Z(n8780) );
  XNOR U8585 ( .A(n8779), .B(n8783), .Z(n8781) );
  XOR U8586 ( .A(n8557), .B(n8784), .Z(n8551) );
  IV U8587 ( .A(n8556), .Z(n8784) );
  XNOR U8588 ( .A(n8553), .B(n8706), .Z(n8556) );
  AND U8589 ( .A(n11049), .B(n5561), .Z(n8706) );
  XOR U8590 ( .A(n8785), .B(n8786), .Z(n8553) );
  ANDN U8591 ( .A(n8787), .B(n8788), .Z(n8786) );
  XNOR U8592 ( .A(n8785), .B(n8789), .Z(n8787) );
  XOR U8593 ( .A(n8563), .B(n8790), .Z(n8557) );
  IV U8594 ( .A(n8562), .Z(n8790) );
  XNOR U8595 ( .A(n8559), .B(n8699), .Z(n8562) );
  AND U8596 ( .A(n11341), .B(n5030), .Z(n8699) );
  XOR U8597 ( .A(n8791), .B(n8792), .Z(n8559) );
  ANDN U8598 ( .A(n8793), .B(n8794), .Z(n8792) );
  XNOR U8599 ( .A(n8791), .B(n8795), .Z(n8793) );
  XOR U8600 ( .A(n8569), .B(n8796), .Z(n8563) );
  IV U8601 ( .A(n8568), .Z(n8796) );
  XNOR U8602 ( .A(n8565), .B(n8692), .Z(n8568) );
  AND U8603 ( .A(n11607), .B(n4525), .Z(n8692) );
  XOR U8604 ( .A(n8797), .B(n8798), .Z(n8565) );
  ANDN U8605 ( .A(n8799), .B(n8800), .Z(n8798) );
  XNOR U8606 ( .A(n8797), .B(n8801), .Z(n8799) );
  XOR U8607 ( .A(n8575), .B(n8802), .Z(n8569) );
  IV U8608 ( .A(n8574), .Z(n8802) );
  XNOR U8609 ( .A(n8571), .B(n8685), .Z(n8574) );
  AND U8610 ( .A(n11869), .B(n4046), .Z(n8685) );
  XOR U8611 ( .A(n8803), .B(n8804), .Z(n8571) );
  ANDN U8612 ( .A(n8805), .B(n8806), .Z(n8804) );
  XNOR U8613 ( .A(n8803), .B(n8807), .Z(n8805) );
  XOR U8614 ( .A(n8581), .B(n8808), .Z(n8575) );
  IV U8615 ( .A(n8580), .Z(n8808) );
  XNOR U8616 ( .A(n8577), .B(n8678), .Z(n8580) );
  AND U8617 ( .A(n12128), .B(n3593), .Z(n8678) );
  XOR U8618 ( .A(n8809), .B(n8810), .Z(n8577) );
  ANDN U8619 ( .A(n8811), .B(n8812), .Z(n8810) );
  XNOR U8620 ( .A(n8809), .B(n8813), .Z(n8811) );
  XOR U8621 ( .A(n8587), .B(n8814), .Z(n8581) );
  IV U8622 ( .A(n8586), .Z(n8814) );
  XNOR U8623 ( .A(n8583), .B(n8671), .Z(n8586) );
  AND U8624 ( .A(n12387), .B(n3166), .Z(n8671) );
  XOR U8625 ( .A(n8815), .B(n8816), .Z(n8583) );
  ANDN U8626 ( .A(n8817), .B(n8818), .Z(n8816) );
  XNOR U8627 ( .A(n8815), .B(n8819), .Z(n8817) );
  XOR U8628 ( .A(n8593), .B(n8820), .Z(n8587) );
  IV U8629 ( .A(n8592), .Z(n8820) );
  XNOR U8630 ( .A(n8589), .B(n8664), .Z(n8592) );
  AND U8631 ( .A(n12644), .B(n2765), .Z(n8664) );
  XOR U8632 ( .A(n8821), .B(n8822), .Z(n8589) );
  ANDN U8633 ( .A(n8823), .B(n8824), .Z(n8822) );
  XNOR U8634 ( .A(n8821), .B(n8825), .Z(n8823) );
  XOR U8635 ( .A(n8599), .B(n8826), .Z(n8593) );
  IV U8636 ( .A(n8598), .Z(n8826) );
  XNOR U8637 ( .A(n8595), .B(n8657), .Z(n8598) );
  AND U8638 ( .A(n12880), .B(n2396), .Z(n8657) );
  XOR U8639 ( .A(n8827), .B(n8828), .Z(n8595) );
  ANDN U8640 ( .A(n8829), .B(n8830), .Z(n8828) );
  XNOR U8641 ( .A(n8827), .B(n8831), .Z(n8829) );
  XOR U8642 ( .A(n8605), .B(n8832), .Z(n8599) );
  IV U8643 ( .A(n8604), .Z(n8832) );
  XNOR U8644 ( .A(n8601), .B(n8650), .Z(n8604) );
  AND U8645 ( .A(n13070), .B(n2053), .Z(n8650) );
  XOR U8646 ( .A(n8833), .B(n8834), .Z(n8601) );
  ANDN U8647 ( .A(n8835), .B(n8836), .Z(n8834) );
  XNOR U8648 ( .A(n8833), .B(n8837), .Z(n8835) );
  XOR U8649 ( .A(n8611), .B(n8838), .Z(n8605) );
  IV U8650 ( .A(n8610), .Z(n8838) );
  XNOR U8651 ( .A(n8607), .B(n8643), .Z(n8610) );
  AND U8652 ( .A(n13207), .B(n1737), .Z(n8643) );
  XOR U8653 ( .A(n8839), .B(n8840), .Z(n8607) );
  ANDN U8654 ( .A(n8841), .B(n8842), .Z(n8840) );
  XNOR U8655 ( .A(n8839), .B(n8843), .Z(n8841) );
  XNOR U8656 ( .A(n8616), .B(n8402), .Z(n8611) );
  XNOR U8657 ( .A(n8613), .B(n8844), .Z(n8616) );
  AND U8658 ( .A(n6527), .B(n1448), .Z(n8844) );
  XOR U8659 ( .A(n8845), .B(n8846), .Z(n8613) );
  ANDN U8660 ( .A(n8847), .B(n8848), .Z(n8846) );
  XNOR U8661 ( .A(n8640), .B(n8845), .Z(n8847) );
  XOR U8662 ( .A(n8849), .B(n8402), .Z(n8637) );
  NANDN U8663 ( .B(n6808), .A(n1185), .Z(n8402) );
  XOR U8664 ( .A(n8850), .B(n8851), .Z(n1185) );
  AND U8665 ( .A(n6809), .B(n8852), .Z(n8851) );
  XNOR U8666 ( .A(n8850), .B(n8623), .Z(n8852) );
  XOR U8667 ( .A(n8621), .B(n8850), .Z(n8623) );
  XOR U8668 ( .A(n8853), .B(n8854), .Z(n8621) );
  ANDN U8669 ( .A(n8853), .B(n8855), .Z(n8854) );
  XOR U8670 ( .A(n8856), .B(n7368), .Z(n8850) );
  IV U8671 ( .A(n8625), .Z(n8849) );
  XOR U8672 ( .A(n8857), .B(n8858), .Z(n8625) );
  AND U8673 ( .A(n8859), .B(n8860), .Z(n8858) );
  XOR U8674 ( .A(n8861), .B(n8857), .Z(n8860) );
  XOR U8675 ( .A(n8629), .B(n8633), .Z(n8636) );
  XOR U8676 ( .A(n8862), .B(n8863), .Z(n8629) );
  IV U8677 ( .A(n8864), .Z(n8863) );
  XOR U8678 ( .A(n8865), .B(n8866), .Z(n8633) );
  AND U8679 ( .A(n8865), .B(n8867), .Z(n8866) );
  XOR U8680 ( .A(n8868), .B(n8859), .Z(n8867) );
  XOR U8681 ( .A(n8869), .B(n8641), .Z(n8859) );
  XOR U8682 ( .A(n8648), .B(n8870), .Z(n8641) );
  IV U8683 ( .A(n8646), .Z(n8870) );
  XNOR U8684 ( .A(n8871), .B(n8645), .Z(n8646) );
  OR U8685 ( .A(n8872), .B(n8873), .Z(n8645) );
  NANDN U8686 ( .B(n6541), .A(n1737), .Z(n8871) );
  XOR U8687 ( .A(n8655), .B(n8874), .Z(n8648) );
  IV U8688 ( .A(n8654), .Z(n8874) );
  XNOR U8689 ( .A(n8651), .B(n8875), .Z(n8654) );
  XOR U8690 ( .A(n8876), .B(n8877), .Z(n8651) );
  NANDN U8691 ( .B(n8878), .A(n8879), .Z(n8876) );
  XOR U8692 ( .A(n8877), .B(n8880), .Z(n8879) );
  XOR U8693 ( .A(n8662), .B(n8881), .Z(n8655) );
  IV U8694 ( .A(n8661), .Z(n8881) );
  XNOR U8695 ( .A(n8658), .B(n8882), .Z(n8661) );
  XOR U8696 ( .A(n8883), .B(n8884), .Z(n8658) );
  ANDN U8697 ( .A(n8885), .B(n8886), .Z(n8884) );
  XNOR U8698 ( .A(n8883), .B(n8887), .Z(n8885) );
  XOR U8699 ( .A(n8669), .B(n8888), .Z(n8662) );
  IV U8700 ( .A(n8668), .Z(n8888) );
  XNOR U8701 ( .A(n8665), .B(n8889), .Z(n8668) );
  XOR U8702 ( .A(n8890), .B(n8891), .Z(n8665) );
  ANDN U8703 ( .A(n8892), .B(n8893), .Z(n8891) );
  XNOR U8704 ( .A(n8890), .B(n8894), .Z(n8892) );
  XOR U8705 ( .A(n8676), .B(n8895), .Z(n8669) );
  IV U8706 ( .A(n8675), .Z(n8895) );
  XNOR U8707 ( .A(n8672), .B(n8896), .Z(n8675) );
  XOR U8708 ( .A(n8897), .B(n8898), .Z(n8672) );
  ANDN U8709 ( .A(n8899), .B(n8900), .Z(n8898) );
  XNOR U8710 ( .A(n8897), .B(n8901), .Z(n8899) );
  XOR U8711 ( .A(n8683), .B(n8902), .Z(n8676) );
  IV U8712 ( .A(n8682), .Z(n8902) );
  XNOR U8713 ( .A(n8679), .B(n8903), .Z(n8682) );
  XOR U8714 ( .A(n8904), .B(n8905), .Z(n8679) );
  ANDN U8715 ( .A(n8906), .B(n8907), .Z(n8905) );
  XNOR U8716 ( .A(n8904), .B(n8908), .Z(n8906) );
  XOR U8717 ( .A(n8690), .B(n8909), .Z(n8683) );
  IV U8718 ( .A(n8689), .Z(n8909) );
  XNOR U8719 ( .A(n8686), .B(n8910), .Z(n8689) );
  XOR U8720 ( .A(n8911), .B(n8912), .Z(n8686) );
  ANDN U8721 ( .A(n8913), .B(n8914), .Z(n8912) );
  XNOR U8722 ( .A(n8911), .B(n8915), .Z(n8913) );
  XOR U8723 ( .A(n8697), .B(n8916), .Z(n8690) );
  IV U8724 ( .A(n8696), .Z(n8916) );
  XNOR U8725 ( .A(n8693), .B(n8917), .Z(n8696) );
  XOR U8726 ( .A(n8918), .B(n8919), .Z(n8693) );
  ANDN U8727 ( .A(n8920), .B(n8921), .Z(n8919) );
  XNOR U8728 ( .A(n8918), .B(n8922), .Z(n8920) );
  XOR U8729 ( .A(n8704), .B(n8923), .Z(n8697) );
  IV U8730 ( .A(n8703), .Z(n8923) );
  XNOR U8731 ( .A(n8700), .B(n8924), .Z(n8703) );
  XOR U8732 ( .A(n8925), .B(n8926), .Z(n8700) );
  ANDN U8733 ( .A(n8927), .B(n8928), .Z(n8926) );
  XNOR U8734 ( .A(n8925), .B(n8929), .Z(n8927) );
  XOR U8735 ( .A(n8711), .B(n8930), .Z(n8704) );
  IV U8736 ( .A(n8710), .Z(n8930) );
  XNOR U8737 ( .A(n8707), .B(n8931), .Z(n8710) );
  XOR U8738 ( .A(n8932), .B(n8933), .Z(n8707) );
  ANDN U8739 ( .A(n8934), .B(n8935), .Z(n8933) );
  XNOR U8740 ( .A(n8932), .B(n8936), .Z(n8934) );
  XOR U8741 ( .A(n8718), .B(n8937), .Z(n8711) );
  IV U8742 ( .A(n8717), .Z(n8937) );
  XNOR U8743 ( .A(n8714), .B(n8938), .Z(n8717) );
  XOR U8744 ( .A(n8939), .B(n8940), .Z(n8714) );
  ANDN U8745 ( .A(n8941), .B(n8942), .Z(n8940) );
  XNOR U8746 ( .A(n8939), .B(n8943), .Z(n8941) );
  XOR U8747 ( .A(n8725), .B(n8944), .Z(n8718) );
  IV U8748 ( .A(n8724), .Z(n8944) );
  XNOR U8749 ( .A(n8721), .B(n8945), .Z(n8724) );
  XOR U8750 ( .A(n8946), .B(n8947), .Z(n8721) );
  ANDN U8751 ( .A(n8948), .B(n8949), .Z(n8947) );
  XNOR U8752 ( .A(n8946), .B(n8950), .Z(n8948) );
  XOR U8753 ( .A(n8732), .B(n8951), .Z(n8725) );
  IV U8754 ( .A(n8731), .Z(n8951) );
  XNOR U8755 ( .A(n8728), .B(n8952), .Z(n8731) );
  XOR U8756 ( .A(n8953), .B(n8954), .Z(n8728) );
  ANDN U8757 ( .A(n8955), .B(n8956), .Z(n8954) );
  XNOR U8758 ( .A(n8953), .B(n8957), .Z(n8955) );
  XOR U8759 ( .A(n8739), .B(n8958), .Z(n8732) );
  IV U8760 ( .A(n8738), .Z(n8958) );
  XNOR U8761 ( .A(n8735), .B(n8959), .Z(n8738) );
  XOR U8762 ( .A(n8960), .B(n8961), .Z(n8735) );
  ANDN U8763 ( .A(n8962), .B(n8963), .Z(n8961) );
  XNOR U8764 ( .A(n8960), .B(n8964), .Z(n8962) );
  XOR U8765 ( .A(n8746), .B(n8965), .Z(n8739) );
  IV U8766 ( .A(n8745), .Z(n8965) );
  XNOR U8767 ( .A(n8742), .B(n8966), .Z(n8745) );
  XOR U8768 ( .A(n8967), .B(n8968), .Z(n8742) );
  ANDN U8769 ( .A(n8969), .B(n8970), .Z(n8968) );
  XNOR U8770 ( .A(n8967), .B(n8971), .Z(n8969) );
  XOR U8771 ( .A(n8753), .B(n8972), .Z(n8746) );
  IV U8772 ( .A(n8752), .Z(n8972) );
  XNOR U8773 ( .A(n8749), .B(n8973), .Z(n8752) );
  XOR U8774 ( .A(n8974), .B(n8975), .Z(n8749) );
  ANDN U8775 ( .A(n8976), .B(n8977), .Z(n8975) );
  XNOR U8776 ( .A(n8974), .B(n8978), .Z(n8976) );
  XOR U8777 ( .A(n8759), .B(n8979), .Z(n8753) );
  IV U8778 ( .A(n8758), .Z(n8979) );
  XNOR U8779 ( .A(n8755), .B(n8973), .Z(n8758) );
  AND U8780 ( .A(n9198), .B(n8748), .Z(n8973) );
  XOR U8781 ( .A(n8980), .B(n8981), .Z(n8755) );
  ANDN U8782 ( .A(n8982), .B(n8983), .Z(n8981) );
  XNOR U8783 ( .A(n8980), .B(n8984), .Z(n8982) );
  XOR U8784 ( .A(n8765), .B(n8985), .Z(n8759) );
  IV U8785 ( .A(n8764), .Z(n8985) );
  XNOR U8786 ( .A(n8761), .B(n8966), .Z(n8764) );
  AND U8787 ( .A(n9621), .B(n8272), .Z(n8966) );
  XOR U8788 ( .A(n8986), .B(n8987), .Z(n8761) );
  ANDN U8789 ( .A(n8988), .B(n8989), .Z(n8987) );
  XNOR U8790 ( .A(n8986), .B(n8990), .Z(n8988) );
  XOR U8791 ( .A(n8771), .B(n8991), .Z(n8765) );
  IV U8792 ( .A(n8770), .Z(n8991) );
  XNOR U8793 ( .A(n8767), .B(n8959), .Z(n8770) );
  AND U8794 ( .A(n10017), .B(n7770), .Z(n8959) );
  XOR U8795 ( .A(n8992), .B(n8993), .Z(n8767) );
  ANDN U8796 ( .A(n8994), .B(n8995), .Z(n8993) );
  XNOR U8797 ( .A(n8992), .B(n8996), .Z(n8994) );
  XOR U8798 ( .A(n8777), .B(n8997), .Z(n8771) );
  IV U8799 ( .A(n8776), .Z(n8997) );
  XNOR U8800 ( .A(n8773), .B(n8952), .Z(n8776) );
  AND U8801 ( .A(n10387), .B(n7241), .Z(n8952) );
  XOR U8802 ( .A(n8998), .B(n8999), .Z(n8773) );
  ANDN U8803 ( .A(n9000), .B(n9001), .Z(n8999) );
  XNOR U8804 ( .A(n8998), .B(n9002), .Z(n9000) );
  XOR U8805 ( .A(n8783), .B(n9003), .Z(n8777) );
  IV U8806 ( .A(n8782), .Z(n9003) );
  XNOR U8807 ( .A(n8779), .B(n8945), .Z(n8782) );
  AND U8808 ( .A(n10731), .B(n6688), .Z(n8945) );
  XOR U8809 ( .A(n9004), .B(n9005), .Z(n8779) );
  ANDN U8810 ( .A(n9006), .B(n9007), .Z(n9005) );
  XNOR U8811 ( .A(n9004), .B(n9008), .Z(n9006) );
  XOR U8812 ( .A(n8789), .B(n9009), .Z(n8783) );
  IV U8813 ( .A(n8788), .Z(n9009) );
  XNOR U8814 ( .A(n8785), .B(n8938), .Z(n8788) );
  AND U8815 ( .A(n11049), .B(n6118), .Z(n8938) );
  XOR U8816 ( .A(n9010), .B(n9011), .Z(n8785) );
  ANDN U8817 ( .A(n9012), .B(n9013), .Z(n9011) );
  XNOR U8818 ( .A(n9010), .B(n9014), .Z(n9012) );
  XOR U8819 ( .A(n8795), .B(n9015), .Z(n8789) );
  IV U8820 ( .A(n8794), .Z(n9015) );
  XNOR U8821 ( .A(n8791), .B(n8931), .Z(n8794) );
  AND U8822 ( .A(n11341), .B(n5561), .Z(n8931) );
  XOR U8823 ( .A(n9016), .B(n9017), .Z(n8791) );
  ANDN U8824 ( .A(n9018), .B(n9019), .Z(n9017) );
  XNOR U8825 ( .A(n9016), .B(n9020), .Z(n9018) );
  XOR U8826 ( .A(n8801), .B(n9021), .Z(n8795) );
  IV U8827 ( .A(n8800), .Z(n9021) );
  XNOR U8828 ( .A(n8797), .B(n8924), .Z(n8800) );
  AND U8829 ( .A(n11607), .B(n5030), .Z(n8924) );
  XOR U8830 ( .A(n9022), .B(n9023), .Z(n8797) );
  ANDN U8831 ( .A(n9024), .B(n9025), .Z(n9023) );
  XNOR U8832 ( .A(n9022), .B(n9026), .Z(n9024) );
  XOR U8833 ( .A(n8807), .B(n9027), .Z(n8801) );
  IV U8834 ( .A(n8806), .Z(n9027) );
  XNOR U8835 ( .A(n8803), .B(n8917), .Z(n8806) );
  AND U8836 ( .A(n11869), .B(n4525), .Z(n8917) );
  XOR U8837 ( .A(n9028), .B(n9029), .Z(n8803) );
  ANDN U8838 ( .A(n9030), .B(n9031), .Z(n9029) );
  XNOR U8839 ( .A(n9028), .B(n9032), .Z(n9030) );
  XOR U8840 ( .A(n8813), .B(n9033), .Z(n8807) );
  IV U8841 ( .A(n8812), .Z(n9033) );
  XNOR U8842 ( .A(n8809), .B(n8910), .Z(n8812) );
  AND U8843 ( .A(n12128), .B(n4046), .Z(n8910) );
  XOR U8844 ( .A(n9034), .B(n9035), .Z(n8809) );
  ANDN U8845 ( .A(n9036), .B(n9037), .Z(n9035) );
  XNOR U8846 ( .A(n9034), .B(n9038), .Z(n9036) );
  XOR U8847 ( .A(n8819), .B(n9039), .Z(n8813) );
  IV U8848 ( .A(n8818), .Z(n9039) );
  XNOR U8849 ( .A(n8815), .B(n8903), .Z(n8818) );
  AND U8850 ( .A(n12387), .B(n3593), .Z(n8903) );
  XOR U8851 ( .A(n9040), .B(n9041), .Z(n8815) );
  ANDN U8852 ( .A(n9042), .B(n9043), .Z(n9041) );
  XNOR U8853 ( .A(n9040), .B(n9044), .Z(n9042) );
  XOR U8854 ( .A(n8825), .B(n9045), .Z(n8819) );
  IV U8855 ( .A(n8824), .Z(n9045) );
  XNOR U8856 ( .A(n8821), .B(n8896), .Z(n8824) );
  AND U8857 ( .A(n12644), .B(n3166), .Z(n8896) );
  XOR U8858 ( .A(n9046), .B(n9047), .Z(n8821) );
  ANDN U8859 ( .A(n9048), .B(n9049), .Z(n9047) );
  XNOR U8860 ( .A(n9046), .B(n9050), .Z(n9048) );
  XOR U8861 ( .A(n8831), .B(n9051), .Z(n8825) );
  IV U8862 ( .A(n8830), .Z(n9051) );
  XNOR U8863 ( .A(n8827), .B(n8889), .Z(n8830) );
  AND U8864 ( .A(n12880), .B(n2765), .Z(n8889) );
  XOR U8865 ( .A(n9052), .B(n9053), .Z(n8827) );
  ANDN U8866 ( .A(n9054), .B(n9055), .Z(n9053) );
  XNOR U8867 ( .A(n9052), .B(n9056), .Z(n9054) );
  XOR U8868 ( .A(n8837), .B(n9057), .Z(n8831) );
  IV U8869 ( .A(n8836), .Z(n9057) );
  XNOR U8870 ( .A(n8833), .B(n8882), .Z(n8836) );
  AND U8871 ( .A(n13070), .B(n2396), .Z(n8882) );
  XOR U8872 ( .A(n9058), .B(n9059), .Z(n8833) );
  ANDN U8873 ( .A(n9060), .B(n9061), .Z(n9059) );
  XNOR U8874 ( .A(n9058), .B(n9062), .Z(n9060) );
  XOR U8875 ( .A(n8843), .B(n9063), .Z(n8837) );
  IV U8876 ( .A(n8842), .Z(n9063) );
  XNOR U8877 ( .A(n8839), .B(n8875), .Z(n8842) );
  AND U8878 ( .A(n13207), .B(n2053), .Z(n8875) );
  XOR U8879 ( .A(n9064), .B(n9065), .Z(n8839) );
  ANDN U8880 ( .A(n9066), .B(n9067), .Z(n9065) );
  XNOR U8881 ( .A(n9064), .B(n9068), .Z(n9066) );
  XNOR U8882 ( .A(n8848), .B(n8640), .Z(n8843) );
  XNOR U8883 ( .A(n8845), .B(n9069), .Z(n8848) );
  AND U8884 ( .A(n6527), .B(n1737), .Z(n9069) );
  XOR U8885 ( .A(n9070), .B(n9071), .Z(n8845) );
  ANDN U8886 ( .A(n9072), .B(n9073), .Z(n9071) );
  XNOR U8887 ( .A(n8872), .B(n9070), .Z(n9072) );
  XOR U8888 ( .A(n9074), .B(n8640), .Z(n8869) );
  NANDN U8889 ( .B(n6808), .A(n1448), .Z(n8640) );
  XOR U8890 ( .A(n9075), .B(n9076), .Z(n1448) );
  AND U8891 ( .A(n6809), .B(n9077), .Z(n9076) );
  XNOR U8892 ( .A(n9075), .B(n8855), .Z(n9077) );
  XOR U8893 ( .A(n8853), .B(n9075), .Z(n8855) );
  XOR U8894 ( .A(n9078), .B(n9079), .Z(n8853) );
  ANDN U8895 ( .A(n9078), .B(n9080), .Z(n9079) );
  XOR U8896 ( .A(n9081), .B(n7368), .Z(n9075) );
  IV U8897 ( .A(n8857), .Z(n9074) );
  XOR U8898 ( .A(n9082), .B(n9083), .Z(n8857) );
  AND U8899 ( .A(n9084), .B(n9085), .Z(n9083) );
  XOR U8900 ( .A(n9086), .B(n9082), .Z(n9085) );
  XOR U8901 ( .A(n8861), .B(n8865), .Z(n8868) );
  XOR U8902 ( .A(n9087), .B(n9088), .Z(n8861) );
  IV U8903 ( .A(n9089), .Z(n9088) );
  XOR U8904 ( .A(n9090), .B(n9091), .Z(n8865) );
  AND U8905 ( .A(n9090), .B(n9092), .Z(n9091) );
  XOR U8906 ( .A(n9093), .B(n9084), .Z(n9092) );
  XOR U8907 ( .A(n9094), .B(n8873), .Z(n9084) );
  XOR U8908 ( .A(n8880), .B(n9095), .Z(n8873) );
  IV U8909 ( .A(n8878), .Z(n9095) );
  XNOR U8910 ( .A(n9096), .B(n8877), .Z(n8878) );
  OR U8911 ( .A(n9097), .B(n9098), .Z(n8877) );
  NANDN U8912 ( .B(n6541), .A(n2053), .Z(n9096) );
  XOR U8913 ( .A(n8887), .B(n9099), .Z(n8880) );
  IV U8914 ( .A(n8886), .Z(n9099) );
  XNOR U8915 ( .A(n8883), .B(n9100), .Z(n8886) );
  XOR U8916 ( .A(n9101), .B(n9102), .Z(n8883) );
  NANDN U8917 ( .B(n9103), .A(n9104), .Z(n9101) );
  XOR U8918 ( .A(n9102), .B(n9105), .Z(n9104) );
  XOR U8919 ( .A(n8894), .B(n9106), .Z(n8887) );
  IV U8920 ( .A(n8893), .Z(n9106) );
  XNOR U8921 ( .A(n8890), .B(n9107), .Z(n8893) );
  XOR U8922 ( .A(n9108), .B(n9109), .Z(n8890) );
  ANDN U8923 ( .A(n9110), .B(n9111), .Z(n9109) );
  XNOR U8924 ( .A(n9108), .B(n9112), .Z(n9110) );
  XOR U8925 ( .A(n8901), .B(n9113), .Z(n8894) );
  IV U8926 ( .A(n8900), .Z(n9113) );
  XNOR U8927 ( .A(n8897), .B(n9114), .Z(n8900) );
  XOR U8928 ( .A(n9115), .B(n9116), .Z(n8897) );
  ANDN U8929 ( .A(n9117), .B(n9118), .Z(n9116) );
  XNOR U8930 ( .A(n9115), .B(n9119), .Z(n9117) );
  XOR U8931 ( .A(n8908), .B(n9120), .Z(n8901) );
  IV U8932 ( .A(n8907), .Z(n9120) );
  XNOR U8933 ( .A(n8904), .B(n9121), .Z(n8907) );
  XOR U8934 ( .A(n9122), .B(n9123), .Z(n8904) );
  ANDN U8935 ( .A(n9124), .B(n9125), .Z(n9123) );
  XNOR U8936 ( .A(n9122), .B(n9126), .Z(n9124) );
  XOR U8937 ( .A(n8915), .B(n9127), .Z(n8908) );
  IV U8938 ( .A(n8914), .Z(n9127) );
  XNOR U8939 ( .A(n8911), .B(n9128), .Z(n8914) );
  XOR U8940 ( .A(n9129), .B(n9130), .Z(n8911) );
  ANDN U8941 ( .A(n9131), .B(n9132), .Z(n9130) );
  XNOR U8942 ( .A(n9129), .B(n9133), .Z(n9131) );
  XOR U8943 ( .A(n8922), .B(n9134), .Z(n8915) );
  IV U8944 ( .A(n8921), .Z(n9134) );
  XNOR U8945 ( .A(n8918), .B(n9135), .Z(n8921) );
  XOR U8946 ( .A(n9136), .B(n9137), .Z(n8918) );
  ANDN U8947 ( .A(n9138), .B(n9139), .Z(n9137) );
  XNOR U8948 ( .A(n9136), .B(n9140), .Z(n9138) );
  XOR U8949 ( .A(n8929), .B(n9141), .Z(n8922) );
  IV U8950 ( .A(n8928), .Z(n9141) );
  XNOR U8951 ( .A(n8925), .B(n9142), .Z(n8928) );
  XOR U8952 ( .A(n9143), .B(n9144), .Z(n8925) );
  ANDN U8953 ( .A(n9145), .B(n9146), .Z(n9144) );
  XNOR U8954 ( .A(n9143), .B(n9147), .Z(n9145) );
  XOR U8955 ( .A(n8936), .B(n9148), .Z(n8929) );
  IV U8956 ( .A(n8935), .Z(n9148) );
  XNOR U8957 ( .A(n8932), .B(n9149), .Z(n8935) );
  XOR U8958 ( .A(n9150), .B(n9151), .Z(n8932) );
  ANDN U8959 ( .A(n9152), .B(n9153), .Z(n9151) );
  XNOR U8960 ( .A(n9150), .B(n9154), .Z(n9152) );
  XOR U8961 ( .A(n8943), .B(n9155), .Z(n8936) );
  IV U8962 ( .A(n8942), .Z(n9155) );
  XNOR U8963 ( .A(n8939), .B(n9156), .Z(n8942) );
  XOR U8964 ( .A(n9157), .B(n9158), .Z(n8939) );
  ANDN U8965 ( .A(n9159), .B(n9160), .Z(n9158) );
  XNOR U8966 ( .A(n9157), .B(n9161), .Z(n9159) );
  XOR U8967 ( .A(n8950), .B(n9162), .Z(n8943) );
  IV U8968 ( .A(n8949), .Z(n9162) );
  XNOR U8969 ( .A(n8946), .B(n9163), .Z(n8949) );
  XOR U8970 ( .A(n9164), .B(n9165), .Z(n8946) );
  ANDN U8971 ( .A(n9166), .B(n9167), .Z(n9165) );
  XNOR U8972 ( .A(n9164), .B(n9168), .Z(n9166) );
  XOR U8973 ( .A(n8957), .B(n9169), .Z(n8950) );
  IV U8974 ( .A(n8956), .Z(n9169) );
  XNOR U8975 ( .A(n8953), .B(n9170), .Z(n8956) );
  XOR U8976 ( .A(n9171), .B(n9172), .Z(n8953) );
  ANDN U8977 ( .A(n9173), .B(n9174), .Z(n9172) );
  XNOR U8978 ( .A(n9171), .B(n9175), .Z(n9173) );
  XOR U8979 ( .A(n8964), .B(n9176), .Z(n8957) );
  IV U8980 ( .A(n8963), .Z(n9176) );
  XNOR U8981 ( .A(n8960), .B(n9177), .Z(n8963) );
  XOR U8982 ( .A(n9178), .B(n9179), .Z(n8960) );
  ANDN U8983 ( .A(n9180), .B(n9181), .Z(n9179) );
  XNOR U8984 ( .A(n9178), .B(n9182), .Z(n9180) );
  XOR U8985 ( .A(n8971), .B(n9183), .Z(n8964) );
  IV U8986 ( .A(n8970), .Z(n9183) );
  XNOR U8987 ( .A(n8967), .B(n9184), .Z(n8970) );
  XOR U8988 ( .A(n9185), .B(n9186), .Z(n8967) );
  ANDN U8989 ( .A(n9187), .B(n9188), .Z(n9186) );
  XNOR U8990 ( .A(n9185), .B(n9189), .Z(n9187) );
  XOR U8991 ( .A(n8978), .B(n9190), .Z(n8971) );
  IV U8992 ( .A(n8977), .Z(n9190) );
  XNOR U8993 ( .A(n8974), .B(n9191), .Z(n8977) );
  XOR U8994 ( .A(n9192), .B(n9193), .Z(n8974) );
  ANDN U8995 ( .A(n9194), .B(n9195), .Z(n9193) );
  XNOR U8996 ( .A(n9192), .B(n9196), .Z(n9194) );
  XOR U8997 ( .A(n8984), .B(n9197), .Z(n8978) );
  IV U8998 ( .A(n8983), .Z(n9197) );
  XNOR U8999 ( .A(n8980), .B(n9198), .Z(n8983) );
  XOR U9000 ( .A(n9199), .B(n9200), .Z(n8980) );
  ANDN U9001 ( .A(n9201), .B(n9202), .Z(n9200) );
  XNOR U9002 ( .A(n9199), .B(n9203), .Z(n9201) );
  XOR U9003 ( .A(n8990), .B(n9204), .Z(n8984) );
  IV U9004 ( .A(n8989), .Z(n9204) );
  XNOR U9005 ( .A(n8986), .B(n9191), .Z(n8989) );
  AND U9006 ( .A(n9621), .B(n8748), .Z(n9191) );
  XOR U9007 ( .A(n9205), .B(n9206), .Z(n8986) );
  ANDN U9008 ( .A(n9207), .B(n9208), .Z(n9206) );
  XNOR U9009 ( .A(n9205), .B(n9209), .Z(n9207) );
  XOR U9010 ( .A(n8996), .B(n9210), .Z(n8990) );
  IV U9011 ( .A(n8995), .Z(n9210) );
  XNOR U9012 ( .A(n8992), .B(n9184), .Z(n8995) );
  AND U9013 ( .A(n10017), .B(n8272), .Z(n9184) );
  XOR U9014 ( .A(n9211), .B(n9212), .Z(n8992) );
  ANDN U9015 ( .A(n9213), .B(n9214), .Z(n9212) );
  XNOR U9016 ( .A(n9211), .B(n9215), .Z(n9213) );
  XOR U9017 ( .A(n9002), .B(n9216), .Z(n8996) );
  IV U9018 ( .A(n9001), .Z(n9216) );
  XNOR U9019 ( .A(n8998), .B(n9177), .Z(n9001) );
  AND U9020 ( .A(n10387), .B(n7770), .Z(n9177) );
  XOR U9021 ( .A(n9217), .B(n9218), .Z(n8998) );
  ANDN U9022 ( .A(n9219), .B(n9220), .Z(n9218) );
  XNOR U9023 ( .A(n9217), .B(n9221), .Z(n9219) );
  XOR U9024 ( .A(n9008), .B(n9222), .Z(n9002) );
  IV U9025 ( .A(n9007), .Z(n9222) );
  XNOR U9026 ( .A(n9004), .B(n9170), .Z(n9007) );
  AND U9027 ( .A(n10731), .B(n7241), .Z(n9170) );
  XOR U9028 ( .A(n9223), .B(n9224), .Z(n9004) );
  ANDN U9029 ( .A(n9225), .B(n9226), .Z(n9224) );
  XNOR U9030 ( .A(n9223), .B(n9227), .Z(n9225) );
  XOR U9031 ( .A(n9014), .B(n9228), .Z(n9008) );
  IV U9032 ( .A(n9013), .Z(n9228) );
  XNOR U9033 ( .A(n9010), .B(n9163), .Z(n9013) );
  AND U9034 ( .A(n11049), .B(n6688), .Z(n9163) );
  XOR U9035 ( .A(n9229), .B(n9230), .Z(n9010) );
  ANDN U9036 ( .A(n9231), .B(n9232), .Z(n9230) );
  XNOR U9037 ( .A(n9229), .B(n9233), .Z(n9231) );
  XOR U9038 ( .A(n9020), .B(n9234), .Z(n9014) );
  IV U9039 ( .A(n9019), .Z(n9234) );
  XNOR U9040 ( .A(n9016), .B(n9156), .Z(n9019) );
  AND U9041 ( .A(n11341), .B(n6118), .Z(n9156) );
  XOR U9042 ( .A(n9235), .B(n9236), .Z(n9016) );
  ANDN U9043 ( .A(n9237), .B(n9238), .Z(n9236) );
  XNOR U9044 ( .A(n9235), .B(n9239), .Z(n9237) );
  XOR U9045 ( .A(n9026), .B(n9240), .Z(n9020) );
  IV U9046 ( .A(n9025), .Z(n9240) );
  XNOR U9047 ( .A(n9022), .B(n9149), .Z(n9025) );
  AND U9048 ( .A(n11607), .B(n5561), .Z(n9149) );
  XOR U9049 ( .A(n9241), .B(n9242), .Z(n9022) );
  ANDN U9050 ( .A(n9243), .B(n9244), .Z(n9242) );
  XNOR U9051 ( .A(n9241), .B(n9245), .Z(n9243) );
  XOR U9052 ( .A(n9032), .B(n9246), .Z(n9026) );
  IV U9053 ( .A(n9031), .Z(n9246) );
  XNOR U9054 ( .A(n9028), .B(n9142), .Z(n9031) );
  AND U9055 ( .A(n11869), .B(n5030), .Z(n9142) );
  XOR U9056 ( .A(n9247), .B(n9248), .Z(n9028) );
  ANDN U9057 ( .A(n9249), .B(n9250), .Z(n9248) );
  XNOR U9058 ( .A(n9247), .B(n9251), .Z(n9249) );
  XOR U9059 ( .A(n9038), .B(n9252), .Z(n9032) );
  IV U9060 ( .A(n9037), .Z(n9252) );
  XNOR U9061 ( .A(n9034), .B(n9135), .Z(n9037) );
  AND U9062 ( .A(n12128), .B(n4525), .Z(n9135) );
  XOR U9063 ( .A(n9253), .B(n9254), .Z(n9034) );
  ANDN U9064 ( .A(n9255), .B(n9256), .Z(n9254) );
  XNOR U9065 ( .A(n9253), .B(n9257), .Z(n9255) );
  XOR U9066 ( .A(n9044), .B(n9258), .Z(n9038) );
  IV U9067 ( .A(n9043), .Z(n9258) );
  XNOR U9068 ( .A(n9040), .B(n9128), .Z(n9043) );
  AND U9069 ( .A(n12387), .B(n4046), .Z(n9128) );
  XOR U9070 ( .A(n9259), .B(n9260), .Z(n9040) );
  ANDN U9071 ( .A(n9261), .B(n9262), .Z(n9260) );
  XNOR U9072 ( .A(n9259), .B(n9263), .Z(n9261) );
  XOR U9073 ( .A(n9050), .B(n9264), .Z(n9044) );
  IV U9074 ( .A(n9049), .Z(n9264) );
  XNOR U9075 ( .A(n9046), .B(n9121), .Z(n9049) );
  AND U9076 ( .A(n12644), .B(n3593), .Z(n9121) );
  XOR U9077 ( .A(n9265), .B(n9266), .Z(n9046) );
  ANDN U9078 ( .A(n9267), .B(n9268), .Z(n9266) );
  XNOR U9079 ( .A(n9265), .B(n9269), .Z(n9267) );
  XOR U9080 ( .A(n9056), .B(n9270), .Z(n9050) );
  IV U9081 ( .A(n9055), .Z(n9270) );
  XNOR U9082 ( .A(n9052), .B(n9114), .Z(n9055) );
  AND U9083 ( .A(n12880), .B(n3166), .Z(n9114) );
  XOR U9084 ( .A(n9271), .B(n9272), .Z(n9052) );
  ANDN U9085 ( .A(n9273), .B(n9274), .Z(n9272) );
  XNOR U9086 ( .A(n9271), .B(n9275), .Z(n9273) );
  XOR U9087 ( .A(n9062), .B(n9276), .Z(n9056) );
  IV U9088 ( .A(n9061), .Z(n9276) );
  XNOR U9089 ( .A(n9058), .B(n9107), .Z(n9061) );
  AND U9090 ( .A(n13070), .B(n2765), .Z(n9107) );
  XOR U9091 ( .A(n9277), .B(n9278), .Z(n9058) );
  ANDN U9092 ( .A(n9279), .B(n9280), .Z(n9278) );
  XNOR U9093 ( .A(n9277), .B(n9281), .Z(n9279) );
  XOR U9094 ( .A(n9068), .B(n9282), .Z(n9062) );
  IV U9095 ( .A(n9067), .Z(n9282) );
  XNOR U9096 ( .A(n9064), .B(n9100), .Z(n9067) );
  AND U9097 ( .A(n13207), .B(n2396), .Z(n9100) );
  XOR U9098 ( .A(n9283), .B(n9284), .Z(n9064) );
  ANDN U9099 ( .A(n9285), .B(n9286), .Z(n9284) );
  XNOR U9100 ( .A(n9283), .B(n9287), .Z(n9285) );
  XNOR U9101 ( .A(n9073), .B(n8872), .Z(n9068) );
  XNOR U9102 ( .A(n9070), .B(n9288), .Z(n9073) );
  AND U9103 ( .A(n6527), .B(n2053), .Z(n9288) );
  XOR U9104 ( .A(n9289), .B(n9290), .Z(n9070) );
  ANDN U9105 ( .A(n9291), .B(n9292), .Z(n9290) );
  XNOR U9106 ( .A(n9097), .B(n9289), .Z(n9291) );
  XOR U9107 ( .A(n9293), .B(n8872), .Z(n9094) );
  NANDN U9108 ( .B(n6808), .A(n1737), .Z(n8872) );
  XOR U9109 ( .A(n9294), .B(n9295), .Z(n1737) );
  AND U9110 ( .A(n6809), .B(n9296), .Z(n9295) );
  XNOR U9111 ( .A(n9294), .B(n9080), .Z(n9296) );
  XOR U9112 ( .A(n9078), .B(n9294), .Z(n9080) );
  XOR U9113 ( .A(n9297), .B(n9298), .Z(n9078) );
  ANDN U9114 ( .A(n9297), .B(n9299), .Z(n9298) );
  XOR U9115 ( .A(n9300), .B(n7368), .Z(n9294) );
  IV U9116 ( .A(n9082), .Z(n9293) );
  XOR U9117 ( .A(n9301), .B(n9302), .Z(n9082) );
  AND U9118 ( .A(n9303), .B(n9304), .Z(n9302) );
  XNOR U9119 ( .A(n9305), .B(n9301), .Z(n9304) );
  XOR U9120 ( .A(n9086), .B(n9090), .Z(n9093) );
  XOR U9121 ( .A(n9306), .B(n9307), .Z(n9086) );
  IV U9122 ( .A(n9308), .Z(n9307) );
  XOR U9123 ( .A(n9309), .B(n9310), .Z(n9090) );
  AND U9124 ( .A(n9309), .B(n9311), .Z(n9310) );
  XOR U9125 ( .A(n9312), .B(n9303), .Z(n9311) );
  XOR U9126 ( .A(n9313), .B(n9098), .Z(n9303) );
  XOR U9127 ( .A(n9105), .B(n9314), .Z(n9098) );
  IV U9128 ( .A(n9103), .Z(n9314) );
  XNOR U9129 ( .A(n9315), .B(n9102), .Z(n9103) );
  OR U9130 ( .A(n9316), .B(n9317), .Z(n9102) );
  NANDN U9131 ( .B(n6541), .A(n2396), .Z(n9315) );
  XOR U9132 ( .A(n9112), .B(n9318), .Z(n9105) );
  IV U9133 ( .A(n9111), .Z(n9318) );
  XNOR U9134 ( .A(n9108), .B(n9319), .Z(n9111) );
  XOR U9135 ( .A(n9320), .B(n9321), .Z(n9108) );
  NANDN U9136 ( .B(n9322), .A(n9323), .Z(n9320) );
  XOR U9137 ( .A(n9321), .B(n9324), .Z(n9323) );
  XOR U9138 ( .A(n9119), .B(n9325), .Z(n9112) );
  IV U9139 ( .A(n9118), .Z(n9325) );
  XNOR U9140 ( .A(n9115), .B(n9326), .Z(n9118) );
  XOR U9141 ( .A(n9327), .B(n9328), .Z(n9115) );
  ANDN U9142 ( .A(n9329), .B(n9330), .Z(n9328) );
  XNOR U9143 ( .A(n9327), .B(n9331), .Z(n9329) );
  XOR U9144 ( .A(n9126), .B(n9332), .Z(n9119) );
  IV U9145 ( .A(n9125), .Z(n9332) );
  XNOR U9146 ( .A(n9122), .B(n9333), .Z(n9125) );
  XOR U9147 ( .A(n9334), .B(n9335), .Z(n9122) );
  ANDN U9148 ( .A(n9336), .B(n9337), .Z(n9335) );
  XNOR U9149 ( .A(n9334), .B(n9338), .Z(n9336) );
  XOR U9150 ( .A(n9133), .B(n9339), .Z(n9126) );
  IV U9151 ( .A(n9132), .Z(n9339) );
  XNOR U9152 ( .A(n9129), .B(n9340), .Z(n9132) );
  XOR U9153 ( .A(n9341), .B(n9342), .Z(n9129) );
  ANDN U9154 ( .A(n9343), .B(n9344), .Z(n9342) );
  XNOR U9155 ( .A(n9341), .B(n9345), .Z(n9343) );
  XOR U9156 ( .A(n9140), .B(n9346), .Z(n9133) );
  IV U9157 ( .A(n9139), .Z(n9346) );
  XNOR U9158 ( .A(n9136), .B(n9347), .Z(n9139) );
  XOR U9159 ( .A(n9348), .B(n9349), .Z(n9136) );
  ANDN U9160 ( .A(n9350), .B(n9351), .Z(n9349) );
  XNOR U9161 ( .A(n9348), .B(n9352), .Z(n9350) );
  XOR U9162 ( .A(n9147), .B(n9353), .Z(n9140) );
  IV U9163 ( .A(n9146), .Z(n9353) );
  XNOR U9164 ( .A(n9143), .B(n9354), .Z(n9146) );
  XOR U9165 ( .A(n9355), .B(n9356), .Z(n9143) );
  ANDN U9166 ( .A(n9357), .B(n9358), .Z(n9356) );
  XNOR U9167 ( .A(n9355), .B(n9359), .Z(n9357) );
  XOR U9168 ( .A(n9154), .B(n9360), .Z(n9147) );
  IV U9169 ( .A(n9153), .Z(n9360) );
  XNOR U9170 ( .A(n9150), .B(n9361), .Z(n9153) );
  XOR U9171 ( .A(n9362), .B(n9363), .Z(n9150) );
  ANDN U9172 ( .A(n9364), .B(n9365), .Z(n9363) );
  XNOR U9173 ( .A(n9362), .B(n9366), .Z(n9364) );
  XOR U9174 ( .A(n9161), .B(n9367), .Z(n9154) );
  IV U9175 ( .A(n9160), .Z(n9367) );
  XNOR U9176 ( .A(n9157), .B(n9368), .Z(n9160) );
  XOR U9177 ( .A(n9369), .B(n9370), .Z(n9157) );
  ANDN U9178 ( .A(n9371), .B(n9372), .Z(n9370) );
  XNOR U9179 ( .A(n9369), .B(n9373), .Z(n9371) );
  XOR U9180 ( .A(n9168), .B(n9374), .Z(n9161) );
  IV U9181 ( .A(n9167), .Z(n9374) );
  XNOR U9182 ( .A(n9164), .B(n9375), .Z(n9167) );
  XOR U9183 ( .A(n9376), .B(n9377), .Z(n9164) );
  ANDN U9184 ( .A(n9378), .B(n9379), .Z(n9377) );
  XNOR U9185 ( .A(n9376), .B(n9380), .Z(n9378) );
  XOR U9186 ( .A(n9175), .B(n9381), .Z(n9168) );
  IV U9187 ( .A(n9174), .Z(n9381) );
  XNOR U9188 ( .A(n9171), .B(n9382), .Z(n9174) );
  XOR U9189 ( .A(n9383), .B(n9384), .Z(n9171) );
  ANDN U9190 ( .A(n9385), .B(n9386), .Z(n9384) );
  XNOR U9191 ( .A(n9383), .B(n9387), .Z(n9385) );
  XOR U9192 ( .A(n9182), .B(n9388), .Z(n9175) );
  IV U9193 ( .A(n9181), .Z(n9388) );
  XNOR U9194 ( .A(n9178), .B(n9389), .Z(n9181) );
  XOR U9195 ( .A(n9390), .B(n9391), .Z(n9178) );
  ANDN U9196 ( .A(n9392), .B(n9393), .Z(n9391) );
  XNOR U9197 ( .A(n9390), .B(n9394), .Z(n9392) );
  XOR U9198 ( .A(n9189), .B(n9395), .Z(n9182) );
  IV U9199 ( .A(n9188), .Z(n9395) );
  XNOR U9200 ( .A(n9185), .B(n9396), .Z(n9188) );
  XOR U9201 ( .A(n9397), .B(n9398), .Z(n9185) );
  ANDN U9202 ( .A(n9399), .B(n9400), .Z(n9398) );
  XNOR U9203 ( .A(n9397), .B(n9401), .Z(n9399) );
  XOR U9204 ( .A(n9196), .B(n9402), .Z(n9189) );
  IV U9205 ( .A(n9195), .Z(n9402) );
  XNOR U9206 ( .A(n9192), .B(n9403), .Z(n9195) );
  XOR U9207 ( .A(n9404), .B(n9405), .Z(n9192) );
  ANDN U9208 ( .A(n9406), .B(n9407), .Z(n9405) );
  XNOR U9209 ( .A(n9404), .B(n9408), .Z(n9406) );
  XOR U9210 ( .A(n9203), .B(n9409), .Z(n9196) );
  IV U9211 ( .A(n9202), .Z(n9409) );
  XNOR U9212 ( .A(n9199), .B(n9410), .Z(n9202) );
  XOR U9213 ( .A(n9411), .B(n9412), .Z(n9199) );
  ANDN U9214 ( .A(n9413), .B(n9414), .Z(n9412) );
  XNOR U9215 ( .A(n9411), .B(n9415), .Z(n9413) );
  XOR U9216 ( .A(n9209), .B(n9416), .Z(n9203) );
  IV U9217 ( .A(n9208), .Z(n9416) );
  XNOR U9218 ( .A(n9205), .B(n9410), .Z(n9208) );
  AND U9219 ( .A(n9621), .B(n9198), .Z(n9410) );
  XOR U9220 ( .A(n9417), .B(n9418), .Z(n9205) );
  ANDN U9221 ( .A(n9419), .B(n9420), .Z(n9418) );
  XNOR U9222 ( .A(n9417), .B(n9421), .Z(n9419) );
  XOR U9223 ( .A(n9215), .B(n9422), .Z(n9209) );
  IV U9224 ( .A(n9214), .Z(n9422) );
  XNOR U9225 ( .A(n9211), .B(n9403), .Z(n9214) );
  AND U9226 ( .A(n10017), .B(n8748), .Z(n9403) );
  XOR U9227 ( .A(n9423), .B(n9424), .Z(n9211) );
  ANDN U9228 ( .A(n9425), .B(n9426), .Z(n9424) );
  XNOR U9229 ( .A(n9423), .B(n9427), .Z(n9425) );
  XOR U9230 ( .A(n9221), .B(n9428), .Z(n9215) );
  IV U9231 ( .A(n9220), .Z(n9428) );
  XNOR U9232 ( .A(n9217), .B(n9396), .Z(n9220) );
  AND U9233 ( .A(n10387), .B(n8272), .Z(n9396) );
  XOR U9234 ( .A(n9429), .B(n9430), .Z(n9217) );
  ANDN U9235 ( .A(n9431), .B(n9432), .Z(n9430) );
  XNOR U9236 ( .A(n9429), .B(n9433), .Z(n9431) );
  XOR U9237 ( .A(n9227), .B(n9434), .Z(n9221) );
  IV U9238 ( .A(n9226), .Z(n9434) );
  XNOR U9239 ( .A(n9223), .B(n9389), .Z(n9226) );
  AND U9240 ( .A(n10731), .B(n7770), .Z(n9389) );
  XOR U9241 ( .A(n9435), .B(n9436), .Z(n9223) );
  ANDN U9242 ( .A(n9437), .B(n9438), .Z(n9436) );
  XNOR U9243 ( .A(n9435), .B(n9439), .Z(n9437) );
  XOR U9244 ( .A(n9233), .B(n9440), .Z(n9227) );
  IV U9245 ( .A(n9232), .Z(n9440) );
  XNOR U9246 ( .A(n9229), .B(n9382), .Z(n9232) );
  AND U9247 ( .A(n11049), .B(n7241), .Z(n9382) );
  XOR U9248 ( .A(n9441), .B(n9442), .Z(n9229) );
  ANDN U9249 ( .A(n9443), .B(n9444), .Z(n9442) );
  XNOR U9250 ( .A(n9441), .B(n9445), .Z(n9443) );
  XOR U9251 ( .A(n9239), .B(n9446), .Z(n9233) );
  IV U9252 ( .A(n9238), .Z(n9446) );
  XNOR U9253 ( .A(n9235), .B(n9375), .Z(n9238) );
  AND U9254 ( .A(n11341), .B(n6688), .Z(n9375) );
  XOR U9255 ( .A(n9447), .B(n9448), .Z(n9235) );
  ANDN U9256 ( .A(n9449), .B(n9450), .Z(n9448) );
  XNOR U9257 ( .A(n9447), .B(n9451), .Z(n9449) );
  XOR U9258 ( .A(n9245), .B(n9452), .Z(n9239) );
  IV U9259 ( .A(n9244), .Z(n9452) );
  XNOR U9260 ( .A(n9241), .B(n9368), .Z(n9244) );
  AND U9261 ( .A(n11607), .B(n6118), .Z(n9368) );
  XOR U9262 ( .A(n9453), .B(n9454), .Z(n9241) );
  ANDN U9263 ( .A(n9455), .B(n9456), .Z(n9454) );
  XNOR U9264 ( .A(n9453), .B(n9457), .Z(n9455) );
  XOR U9265 ( .A(n9251), .B(n9458), .Z(n9245) );
  IV U9266 ( .A(n9250), .Z(n9458) );
  XNOR U9267 ( .A(n9247), .B(n9361), .Z(n9250) );
  AND U9268 ( .A(n11869), .B(n5561), .Z(n9361) );
  XOR U9269 ( .A(n9459), .B(n9460), .Z(n9247) );
  ANDN U9270 ( .A(n9461), .B(n9462), .Z(n9460) );
  XNOR U9271 ( .A(n9459), .B(n9463), .Z(n9461) );
  XOR U9272 ( .A(n9257), .B(n9464), .Z(n9251) );
  IV U9273 ( .A(n9256), .Z(n9464) );
  XNOR U9274 ( .A(n9253), .B(n9354), .Z(n9256) );
  AND U9275 ( .A(n12128), .B(n5030), .Z(n9354) );
  XOR U9276 ( .A(n9465), .B(n9466), .Z(n9253) );
  ANDN U9277 ( .A(n9467), .B(n9468), .Z(n9466) );
  XNOR U9278 ( .A(n9465), .B(n9469), .Z(n9467) );
  XOR U9279 ( .A(n9263), .B(n9470), .Z(n9257) );
  IV U9280 ( .A(n9262), .Z(n9470) );
  XNOR U9281 ( .A(n9259), .B(n9347), .Z(n9262) );
  AND U9282 ( .A(n12387), .B(n4525), .Z(n9347) );
  XOR U9283 ( .A(n9471), .B(n9472), .Z(n9259) );
  ANDN U9284 ( .A(n9473), .B(n9474), .Z(n9472) );
  XNOR U9285 ( .A(n9471), .B(n9475), .Z(n9473) );
  XOR U9286 ( .A(n9269), .B(n9476), .Z(n9263) );
  IV U9287 ( .A(n9268), .Z(n9476) );
  XNOR U9288 ( .A(n9265), .B(n9340), .Z(n9268) );
  AND U9289 ( .A(n12644), .B(n4046), .Z(n9340) );
  XOR U9290 ( .A(n9477), .B(n9478), .Z(n9265) );
  ANDN U9291 ( .A(n9479), .B(n9480), .Z(n9478) );
  XNOR U9292 ( .A(n9477), .B(n9481), .Z(n9479) );
  XOR U9293 ( .A(n9275), .B(n9482), .Z(n9269) );
  IV U9294 ( .A(n9274), .Z(n9482) );
  XNOR U9295 ( .A(n9271), .B(n9333), .Z(n9274) );
  AND U9296 ( .A(n12880), .B(n3593), .Z(n9333) );
  XOR U9297 ( .A(n9483), .B(n9484), .Z(n9271) );
  ANDN U9298 ( .A(n9485), .B(n9486), .Z(n9484) );
  XNOR U9299 ( .A(n9483), .B(n9487), .Z(n9485) );
  XOR U9300 ( .A(n9281), .B(n9488), .Z(n9275) );
  IV U9301 ( .A(n9280), .Z(n9488) );
  XNOR U9302 ( .A(n9277), .B(n9326), .Z(n9280) );
  AND U9303 ( .A(n13070), .B(n3166), .Z(n9326) );
  XOR U9304 ( .A(n9489), .B(n9490), .Z(n9277) );
  ANDN U9305 ( .A(n9491), .B(n9492), .Z(n9490) );
  XNOR U9306 ( .A(n9489), .B(n9493), .Z(n9491) );
  XOR U9307 ( .A(n9287), .B(n9494), .Z(n9281) );
  IV U9308 ( .A(n9286), .Z(n9494) );
  XNOR U9309 ( .A(n9283), .B(n9319), .Z(n9286) );
  AND U9310 ( .A(n13207), .B(n2765), .Z(n9319) );
  XOR U9311 ( .A(n9495), .B(n9496), .Z(n9283) );
  ANDN U9312 ( .A(n9497), .B(n9498), .Z(n9496) );
  XNOR U9313 ( .A(n9495), .B(n9499), .Z(n9497) );
  XNOR U9314 ( .A(n9292), .B(n9097), .Z(n9287) );
  XNOR U9315 ( .A(n9289), .B(n9500), .Z(n9292) );
  AND U9316 ( .A(n6527), .B(n2396), .Z(n9500) );
  XOR U9317 ( .A(n9501), .B(n9502), .Z(n9289) );
  ANDN U9318 ( .A(n9503), .B(n9504), .Z(n9502) );
  XNOR U9319 ( .A(n9316), .B(n9501), .Z(n9503) );
  XOR U9320 ( .A(n9505), .B(n9097), .Z(n9313) );
  NANDN U9321 ( .B(n6808), .A(n2053), .Z(n9097) );
  XOR U9322 ( .A(n9506), .B(n9507), .Z(n2053) );
  AND U9323 ( .A(n6809), .B(n9508), .Z(n9507) );
  XNOR U9324 ( .A(n9506), .B(n9299), .Z(n9508) );
  XOR U9325 ( .A(n9297), .B(n9506), .Z(n9299) );
  XOR U9326 ( .A(n9509), .B(n9510), .Z(n9297) );
  ANDN U9327 ( .A(n9509), .B(n9511), .Z(n9510) );
  XOR U9328 ( .A(n9512), .B(n7368), .Z(n9506) );
  IV U9329 ( .A(n9301), .Z(n9505) );
  XOR U9330 ( .A(n9513), .B(n9514), .Z(n9301) );
  AND U9331 ( .A(n9515), .B(n9516), .Z(n9514) );
  XNOR U9332 ( .A(n9517), .B(n9513), .Z(n9516) );
  XNOR U9333 ( .A(n9305), .B(n9309), .Z(n9312) );
  XOR U9334 ( .A(n9518), .B(n9519), .Z(n9305) );
  XOR U9335 ( .A(n9520), .B(n9521), .Z(n9309) );
  AND U9336 ( .A(n9520), .B(n9522), .Z(n9521) );
  XOR U9337 ( .A(n9523), .B(n9515), .Z(n9522) );
  XOR U9338 ( .A(n9524), .B(n9317), .Z(n9515) );
  XOR U9339 ( .A(n9324), .B(n9525), .Z(n9317) );
  IV U9340 ( .A(n9322), .Z(n9525) );
  XNOR U9341 ( .A(n9526), .B(n9321), .Z(n9322) );
  OR U9342 ( .A(n9527), .B(n9528), .Z(n9321) );
  NANDN U9343 ( .B(n6541), .A(n2765), .Z(n9526) );
  XOR U9344 ( .A(n9331), .B(n9529), .Z(n9324) );
  IV U9345 ( .A(n9330), .Z(n9529) );
  XNOR U9346 ( .A(n9327), .B(n9530), .Z(n9330) );
  XOR U9347 ( .A(n9531), .B(n9532), .Z(n9327) );
  NANDN U9348 ( .B(n9533), .A(n9534), .Z(n9531) );
  XOR U9349 ( .A(n9532), .B(n9535), .Z(n9534) );
  XOR U9350 ( .A(n9338), .B(n9536), .Z(n9331) );
  IV U9351 ( .A(n9337), .Z(n9536) );
  XNOR U9352 ( .A(n9334), .B(n9537), .Z(n9337) );
  XOR U9353 ( .A(n9538), .B(n9539), .Z(n9334) );
  ANDN U9354 ( .A(n9540), .B(n9541), .Z(n9539) );
  XNOR U9355 ( .A(n9538), .B(n9542), .Z(n9540) );
  XOR U9356 ( .A(n9345), .B(n9543), .Z(n9338) );
  IV U9357 ( .A(n9344), .Z(n9543) );
  XNOR U9358 ( .A(n9341), .B(n9544), .Z(n9344) );
  XOR U9359 ( .A(n9545), .B(n9546), .Z(n9341) );
  ANDN U9360 ( .A(n9547), .B(n9548), .Z(n9546) );
  XNOR U9361 ( .A(n9545), .B(n9549), .Z(n9547) );
  XOR U9362 ( .A(n9352), .B(n9550), .Z(n9345) );
  IV U9363 ( .A(n9351), .Z(n9550) );
  XNOR U9364 ( .A(n9348), .B(n9551), .Z(n9351) );
  XOR U9365 ( .A(n9552), .B(n9553), .Z(n9348) );
  ANDN U9366 ( .A(n9554), .B(n9555), .Z(n9553) );
  XNOR U9367 ( .A(n9552), .B(n9556), .Z(n9554) );
  XOR U9368 ( .A(n9359), .B(n9557), .Z(n9352) );
  IV U9369 ( .A(n9358), .Z(n9557) );
  XNOR U9370 ( .A(n9355), .B(n9558), .Z(n9358) );
  XOR U9371 ( .A(n9559), .B(n9560), .Z(n9355) );
  ANDN U9372 ( .A(n9561), .B(n9562), .Z(n9560) );
  XNOR U9373 ( .A(n9559), .B(n9563), .Z(n9561) );
  XOR U9374 ( .A(n9366), .B(n9564), .Z(n9359) );
  IV U9375 ( .A(n9365), .Z(n9564) );
  XNOR U9376 ( .A(n9362), .B(n9565), .Z(n9365) );
  XOR U9377 ( .A(n9566), .B(n9567), .Z(n9362) );
  ANDN U9378 ( .A(n9568), .B(n9569), .Z(n9567) );
  XNOR U9379 ( .A(n9566), .B(n9570), .Z(n9568) );
  XOR U9380 ( .A(n9373), .B(n9571), .Z(n9366) );
  IV U9381 ( .A(n9372), .Z(n9571) );
  XNOR U9382 ( .A(n9369), .B(n9572), .Z(n9372) );
  XOR U9383 ( .A(n9573), .B(n9574), .Z(n9369) );
  ANDN U9384 ( .A(n9575), .B(n9576), .Z(n9574) );
  XNOR U9385 ( .A(n9573), .B(n9577), .Z(n9575) );
  XOR U9386 ( .A(n9380), .B(n9578), .Z(n9373) );
  IV U9387 ( .A(n9379), .Z(n9578) );
  XNOR U9388 ( .A(n9376), .B(n9579), .Z(n9379) );
  XOR U9389 ( .A(n9580), .B(n9581), .Z(n9376) );
  ANDN U9390 ( .A(n9582), .B(n9583), .Z(n9581) );
  XNOR U9391 ( .A(n9580), .B(n9584), .Z(n9582) );
  XOR U9392 ( .A(n9387), .B(n9585), .Z(n9380) );
  IV U9393 ( .A(n9386), .Z(n9585) );
  XNOR U9394 ( .A(n9383), .B(n9586), .Z(n9386) );
  XOR U9395 ( .A(n9587), .B(n9588), .Z(n9383) );
  ANDN U9396 ( .A(n9589), .B(n9590), .Z(n9588) );
  XNOR U9397 ( .A(n9587), .B(n9591), .Z(n9589) );
  XOR U9398 ( .A(n9394), .B(n9592), .Z(n9387) );
  IV U9399 ( .A(n9393), .Z(n9592) );
  XNOR U9400 ( .A(n9390), .B(n9593), .Z(n9393) );
  XOR U9401 ( .A(n9594), .B(n9595), .Z(n9390) );
  ANDN U9402 ( .A(n9596), .B(n9597), .Z(n9595) );
  XNOR U9403 ( .A(n9594), .B(n9598), .Z(n9596) );
  XOR U9404 ( .A(n9401), .B(n9599), .Z(n9394) );
  IV U9405 ( .A(n9400), .Z(n9599) );
  XNOR U9406 ( .A(n9397), .B(n9600), .Z(n9400) );
  XOR U9407 ( .A(n9601), .B(n9602), .Z(n9397) );
  ANDN U9408 ( .A(n9603), .B(n9604), .Z(n9602) );
  XNOR U9409 ( .A(n9601), .B(n9605), .Z(n9603) );
  XOR U9410 ( .A(n9408), .B(n9606), .Z(n9401) );
  IV U9411 ( .A(n9407), .Z(n9606) );
  XNOR U9412 ( .A(n9404), .B(n9607), .Z(n9407) );
  XOR U9413 ( .A(n9608), .B(n9609), .Z(n9404) );
  ANDN U9414 ( .A(n9610), .B(n9611), .Z(n9609) );
  XNOR U9415 ( .A(n9608), .B(n9612), .Z(n9610) );
  XOR U9416 ( .A(n9415), .B(n9613), .Z(n9408) );
  IV U9417 ( .A(n9414), .Z(n9613) );
  XNOR U9418 ( .A(n9411), .B(n9614), .Z(n9414) );
  XOR U9419 ( .A(n9615), .B(n9616), .Z(n9411) );
  ANDN U9420 ( .A(n9617), .B(n9618), .Z(n9616) );
  XNOR U9421 ( .A(n9615), .B(n9619), .Z(n9617) );
  XOR U9422 ( .A(n9421), .B(n9620), .Z(n9415) );
  IV U9423 ( .A(n9420), .Z(n9620) );
  XNOR U9424 ( .A(n9417), .B(n9621), .Z(n9420) );
  XOR U9425 ( .A(n9622), .B(n9623), .Z(n9417) );
  ANDN U9426 ( .A(n9624), .B(n9625), .Z(n9623) );
  XNOR U9427 ( .A(n9622), .B(n9626), .Z(n9624) );
  XOR U9428 ( .A(n9427), .B(n9627), .Z(n9421) );
  IV U9429 ( .A(n9426), .Z(n9627) );
  XNOR U9430 ( .A(n9423), .B(n9614), .Z(n9426) );
  AND U9431 ( .A(n10017), .B(n9198), .Z(n9614) );
  XOR U9432 ( .A(n9628), .B(n9629), .Z(n9423) );
  ANDN U9433 ( .A(n9630), .B(n9631), .Z(n9629) );
  XNOR U9434 ( .A(n9628), .B(n9632), .Z(n9630) );
  XOR U9435 ( .A(n9433), .B(n9633), .Z(n9427) );
  IV U9436 ( .A(n9432), .Z(n9633) );
  XNOR U9437 ( .A(n9429), .B(n9607), .Z(n9432) );
  AND U9438 ( .A(n10387), .B(n8748), .Z(n9607) );
  XOR U9439 ( .A(n9634), .B(n9635), .Z(n9429) );
  ANDN U9440 ( .A(n9636), .B(n9637), .Z(n9635) );
  XNOR U9441 ( .A(n9634), .B(n9638), .Z(n9636) );
  XOR U9442 ( .A(n9439), .B(n9639), .Z(n9433) );
  IV U9443 ( .A(n9438), .Z(n9639) );
  XNOR U9444 ( .A(n9435), .B(n9600), .Z(n9438) );
  AND U9445 ( .A(n10731), .B(n8272), .Z(n9600) );
  XOR U9446 ( .A(n9640), .B(n9641), .Z(n9435) );
  ANDN U9447 ( .A(n9642), .B(n9643), .Z(n9641) );
  XNOR U9448 ( .A(n9640), .B(n9644), .Z(n9642) );
  XOR U9449 ( .A(n9445), .B(n9645), .Z(n9439) );
  IV U9450 ( .A(n9444), .Z(n9645) );
  XNOR U9451 ( .A(n9441), .B(n9593), .Z(n9444) );
  AND U9452 ( .A(n11049), .B(n7770), .Z(n9593) );
  XOR U9453 ( .A(n9646), .B(n9647), .Z(n9441) );
  ANDN U9454 ( .A(n9648), .B(n9649), .Z(n9647) );
  XNOR U9455 ( .A(n9646), .B(n9650), .Z(n9648) );
  XOR U9456 ( .A(n9451), .B(n9651), .Z(n9445) );
  IV U9457 ( .A(n9450), .Z(n9651) );
  XNOR U9458 ( .A(n9447), .B(n9586), .Z(n9450) );
  AND U9459 ( .A(n11341), .B(n7241), .Z(n9586) );
  XOR U9460 ( .A(n9652), .B(n9653), .Z(n9447) );
  ANDN U9461 ( .A(n9654), .B(n9655), .Z(n9653) );
  XNOR U9462 ( .A(n9652), .B(n9656), .Z(n9654) );
  XOR U9463 ( .A(n9457), .B(n9657), .Z(n9451) );
  IV U9464 ( .A(n9456), .Z(n9657) );
  XNOR U9465 ( .A(n9453), .B(n9579), .Z(n9456) );
  AND U9466 ( .A(n11607), .B(n6688), .Z(n9579) );
  XOR U9467 ( .A(n9658), .B(n9659), .Z(n9453) );
  ANDN U9468 ( .A(n9660), .B(n9661), .Z(n9659) );
  XNOR U9469 ( .A(n9658), .B(n9662), .Z(n9660) );
  XOR U9470 ( .A(n9463), .B(n9663), .Z(n9457) );
  IV U9471 ( .A(n9462), .Z(n9663) );
  XNOR U9472 ( .A(n9459), .B(n9572), .Z(n9462) );
  AND U9473 ( .A(n11869), .B(n6118), .Z(n9572) );
  XOR U9474 ( .A(n9664), .B(n9665), .Z(n9459) );
  ANDN U9475 ( .A(n9666), .B(n9667), .Z(n9665) );
  XNOR U9476 ( .A(n9664), .B(n9668), .Z(n9666) );
  XOR U9477 ( .A(n9469), .B(n9669), .Z(n9463) );
  IV U9478 ( .A(n9468), .Z(n9669) );
  XNOR U9479 ( .A(n9465), .B(n9565), .Z(n9468) );
  AND U9480 ( .A(n12128), .B(n5561), .Z(n9565) );
  XOR U9481 ( .A(n9670), .B(n9671), .Z(n9465) );
  ANDN U9482 ( .A(n9672), .B(n9673), .Z(n9671) );
  XNOR U9483 ( .A(n9670), .B(n9674), .Z(n9672) );
  XOR U9484 ( .A(n9475), .B(n9675), .Z(n9469) );
  IV U9485 ( .A(n9474), .Z(n9675) );
  XNOR U9486 ( .A(n9471), .B(n9558), .Z(n9474) );
  AND U9487 ( .A(n12387), .B(n5030), .Z(n9558) );
  XOR U9488 ( .A(n9676), .B(n9677), .Z(n9471) );
  ANDN U9489 ( .A(n9678), .B(n9679), .Z(n9677) );
  XNOR U9490 ( .A(n9676), .B(n9680), .Z(n9678) );
  XOR U9491 ( .A(n9481), .B(n9681), .Z(n9475) );
  IV U9492 ( .A(n9480), .Z(n9681) );
  XNOR U9493 ( .A(n9477), .B(n9551), .Z(n9480) );
  AND U9494 ( .A(n12644), .B(n4525), .Z(n9551) );
  XOR U9495 ( .A(n9682), .B(n9683), .Z(n9477) );
  ANDN U9496 ( .A(n9684), .B(n9685), .Z(n9683) );
  XNOR U9497 ( .A(n9682), .B(n9686), .Z(n9684) );
  XOR U9498 ( .A(n9487), .B(n9687), .Z(n9481) );
  IV U9499 ( .A(n9486), .Z(n9687) );
  XNOR U9500 ( .A(n9483), .B(n9544), .Z(n9486) );
  AND U9501 ( .A(n12880), .B(n4046), .Z(n9544) );
  XOR U9502 ( .A(n9688), .B(n9689), .Z(n9483) );
  ANDN U9503 ( .A(n9690), .B(n9691), .Z(n9689) );
  XNOR U9504 ( .A(n9688), .B(n9692), .Z(n9690) );
  XOR U9505 ( .A(n9493), .B(n9693), .Z(n9487) );
  IV U9506 ( .A(n9492), .Z(n9693) );
  XNOR U9507 ( .A(n9489), .B(n9537), .Z(n9492) );
  AND U9508 ( .A(n13070), .B(n3593), .Z(n9537) );
  XOR U9509 ( .A(n9694), .B(n9695), .Z(n9489) );
  ANDN U9510 ( .A(n9696), .B(n9697), .Z(n9695) );
  XNOR U9511 ( .A(n9694), .B(n9698), .Z(n9696) );
  XOR U9512 ( .A(n9499), .B(n9699), .Z(n9493) );
  IV U9513 ( .A(n9498), .Z(n9699) );
  XNOR U9514 ( .A(n9495), .B(n9530), .Z(n9498) );
  AND U9515 ( .A(n13207), .B(n3166), .Z(n9530) );
  XOR U9516 ( .A(n9700), .B(n9701), .Z(n9495) );
  ANDN U9517 ( .A(n9702), .B(n9703), .Z(n9701) );
  XNOR U9518 ( .A(n9700), .B(n9704), .Z(n9702) );
  XNOR U9519 ( .A(n9504), .B(n9316), .Z(n9499) );
  XNOR U9520 ( .A(n9501), .B(n9705), .Z(n9504) );
  AND U9521 ( .A(n6527), .B(n2765), .Z(n9705) );
  XOR U9522 ( .A(n9706), .B(n9707), .Z(n9501) );
  ANDN U9523 ( .A(n9708), .B(n9709), .Z(n9707) );
  XNOR U9524 ( .A(n9527), .B(n9706), .Z(n9708) );
  XOR U9525 ( .A(n9710), .B(n9316), .Z(n9524) );
  NANDN U9526 ( .B(n6808), .A(n2396), .Z(n9316) );
  XOR U9527 ( .A(n9711), .B(n9712), .Z(n2396) );
  AND U9528 ( .A(n6809), .B(n9713), .Z(n9712) );
  XNOR U9529 ( .A(n9711), .B(n9511), .Z(n9713) );
  XOR U9530 ( .A(n9509), .B(n9711), .Z(n9511) );
  XOR U9531 ( .A(n9714), .B(n9715), .Z(n9509) );
  ANDN U9532 ( .A(n9714), .B(n9716), .Z(n9715) );
  XOR U9533 ( .A(n9717), .B(n7368), .Z(n9711) );
  IV U9534 ( .A(n9513), .Z(n9710) );
  XOR U9535 ( .A(n9718), .B(n9719), .Z(n9513) );
  AND U9536 ( .A(n9720), .B(n9721), .Z(n9719) );
  XNOR U9537 ( .A(n9722), .B(n9718), .Z(n9721) );
  XNOR U9538 ( .A(n9517), .B(n9520), .Z(n9523) );
  XOR U9539 ( .A(n9723), .B(n9724), .Z(n9517) );
  XOR U9540 ( .A(n9725), .B(n9726), .Z(n9520) );
  AND U9541 ( .A(n9725), .B(n9727), .Z(n9726) );
  XOR U9542 ( .A(n9728), .B(n9720), .Z(n9727) );
  XOR U9543 ( .A(n9729), .B(n9528), .Z(n9720) );
  XOR U9544 ( .A(n9535), .B(n9730), .Z(n9528) );
  IV U9545 ( .A(n9533), .Z(n9730) );
  XNOR U9546 ( .A(n9731), .B(n9532), .Z(n9533) );
  OR U9547 ( .A(n9732), .B(n9733), .Z(n9532) );
  NANDN U9548 ( .B(n6541), .A(n3166), .Z(n9731) );
  XOR U9549 ( .A(n9542), .B(n9734), .Z(n9535) );
  IV U9550 ( .A(n9541), .Z(n9734) );
  XNOR U9551 ( .A(n9538), .B(n9735), .Z(n9541) );
  XOR U9552 ( .A(n9736), .B(n9737), .Z(n9538) );
  NANDN U9553 ( .B(n9738), .A(n9739), .Z(n9736) );
  XOR U9554 ( .A(n9737), .B(n9740), .Z(n9739) );
  XOR U9555 ( .A(n9549), .B(n9741), .Z(n9542) );
  IV U9556 ( .A(n9548), .Z(n9741) );
  XNOR U9557 ( .A(n9545), .B(n9742), .Z(n9548) );
  XOR U9558 ( .A(n9743), .B(n9744), .Z(n9545) );
  ANDN U9559 ( .A(n9745), .B(n9746), .Z(n9744) );
  XNOR U9560 ( .A(n9743), .B(n9747), .Z(n9745) );
  XOR U9561 ( .A(n9556), .B(n9748), .Z(n9549) );
  IV U9562 ( .A(n9555), .Z(n9748) );
  XNOR U9563 ( .A(n9552), .B(n9749), .Z(n9555) );
  XOR U9564 ( .A(n9750), .B(n9751), .Z(n9552) );
  ANDN U9565 ( .A(n9752), .B(n9753), .Z(n9751) );
  XNOR U9566 ( .A(n9750), .B(n9754), .Z(n9752) );
  XOR U9567 ( .A(n9563), .B(n9755), .Z(n9556) );
  IV U9568 ( .A(n9562), .Z(n9755) );
  XNOR U9569 ( .A(n9559), .B(n9756), .Z(n9562) );
  XOR U9570 ( .A(n9757), .B(n9758), .Z(n9559) );
  ANDN U9571 ( .A(n9759), .B(n9760), .Z(n9758) );
  XNOR U9572 ( .A(n9757), .B(n9761), .Z(n9759) );
  XOR U9573 ( .A(n9570), .B(n9762), .Z(n9563) );
  IV U9574 ( .A(n9569), .Z(n9762) );
  XNOR U9575 ( .A(n9566), .B(n9763), .Z(n9569) );
  XOR U9576 ( .A(n9764), .B(n9765), .Z(n9566) );
  ANDN U9577 ( .A(n9766), .B(n9767), .Z(n9765) );
  XNOR U9578 ( .A(n9764), .B(n9768), .Z(n9766) );
  XOR U9579 ( .A(n9577), .B(n9769), .Z(n9570) );
  IV U9580 ( .A(n9576), .Z(n9769) );
  XNOR U9581 ( .A(n9573), .B(n9770), .Z(n9576) );
  XOR U9582 ( .A(n9771), .B(n9772), .Z(n9573) );
  ANDN U9583 ( .A(n9773), .B(n9774), .Z(n9772) );
  XNOR U9584 ( .A(n9771), .B(n9775), .Z(n9773) );
  XOR U9585 ( .A(n9584), .B(n9776), .Z(n9577) );
  IV U9586 ( .A(n9583), .Z(n9776) );
  XNOR U9587 ( .A(n9580), .B(n9777), .Z(n9583) );
  XOR U9588 ( .A(n9778), .B(n9779), .Z(n9580) );
  ANDN U9589 ( .A(n9780), .B(n9781), .Z(n9779) );
  XNOR U9590 ( .A(n9778), .B(n9782), .Z(n9780) );
  XOR U9591 ( .A(n9591), .B(n9783), .Z(n9584) );
  IV U9592 ( .A(n9590), .Z(n9783) );
  XNOR U9593 ( .A(n9587), .B(n9784), .Z(n9590) );
  XOR U9594 ( .A(n9785), .B(n9786), .Z(n9587) );
  ANDN U9595 ( .A(n9787), .B(n9788), .Z(n9786) );
  XNOR U9596 ( .A(n9785), .B(n9789), .Z(n9787) );
  XOR U9597 ( .A(n9598), .B(n9790), .Z(n9591) );
  IV U9598 ( .A(n9597), .Z(n9790) );
  XNOR U9599 ( .A(n9594), .B(n9791), .Z(n9597) );
  XOR U9600 ( .A(n9792), .B(n9793), .Z(n9594) );
  ANDN U9601 ( .A(n9794), .B(n9795), .Z(n9793) );
  XNOR U9602 ( .A(n9792), .B(n9796), .Z(n9794) );
  XOR U9603 ( .A(n9605), .B(n9797), .Z(n9598) );
  IV U9604 ( .A(n9604), .Z(n9797) );
  XNOR U9605 ( .A(n9601), .B(n9798), .Z(n9604) );
  XOR U9606 ( .A(n9799), .B(n9800), .Z(n9601) );
  ANDN U9607 ( .A(n9801), .B(n9802), .Z(n9800) );
  XNOR U9608 ( .A(n9799), .B(n9803), .Z(n9801) );
  XOR U9609 ( .A(n9612), .B(n9804), .Z(n9605) );
  IV U9610 ( .A(n9611), .Z(n9804) );
  XNOR U9611 ( .A(n9608), .B(n9805), .Z(n9611) );
  XOR U9612 ( .A(n9806), .B(n9807), .Z(n9608) );
  ANDN U9613 ( .A(n9808), .B(n9809), .Z(n9807) );
  XNOR U9614 ( .A(n9806), .B(n9810), .Z(n9808) );
  XOR U9615 ( .A(n9619), .B(n9811), .Z(n9612) );
  IV U9616 ( .A(n9618), .Z(n9811) );
  XNOR U9617 ( .A(n9615), .B(n9812), .Z(n9618) );
  XOR U9618 ( .A(n9813), .B(n9814), .Z(n9615) );
  ANDN U9619 ( .A(n9815), .B(n9816), .Z(n9814) );
  XNOR U9620 ( .A(n9813), .B(n9817), .Z(n9815) );
  XOR U9621 ( .A(n9626), .B(n9818), .Z(n9619) );
  IV U9622 ( .A(n9625), .Z(n9818) );
  XNOR U9623 ( .A(n9622), .B(n9819), .Z(n9625) );
  XOR U9624 ( .A(n9820), .B(n9821), .Z(n9622) );
  ANDN U9625 ( .A(n9822), .B(n9823), .Z(n9821) );
  XNOR U9626 ( .A(n9820), .B(n9824), .Z(n9822) );
  XOR U9627 ( .A(n9632), .B(n9825), .Z(n9626) );
  IV U9628 ( .A(n9631), .Z(n9825) );
  XNOR U9629 ( .A(n9628), .B(n9819), .Z(n9631) );
  AND U9630 ( .A(n10017), .B(n9621), .Z(n9819) );
  XOR U9631 ( .A(n9826), .B(n9827), .Z(n9628) );
  ANDN U9632 ( .A(n9828), .B(n9829), .Z(n9827) );
  XNOR U9633 ( .A(n9826), .B(n9830), .Z(n9828) );
  XOR U9634 ( .A(n9638), .B(n9831), .Z(n9632) );
  IV U9635 ( .A(n9637), .Z(n9831) );
  XNOR U9636 ( .A(n9634), .B(n9812), .Z(n9637) );
  AND U9637 ( .A(n10387), .B(n9198), .Z(n9812) );
  XOR U9638 ( .A(n9832), .B(n9833), .Z(n9634) );
  ANDN U9639 ( .A(n9834), .B(n9835), .Z(n9833) );
  XNOR U9640 ( .A(n9832), .B(n9836), .Z(n9834) );
  XOR U9641 ( .A(n9644), .B(n9837), .Z(n9638) );
  IV U9642 ( .A(n9643), .Z(n9837) );
  XNOR U9643 ( .A(n9640), .B(n9805), .Z(n9643) );
  AND U9644 ( .A(n10731), .B(n8748), .Z(n9805) );
  XOR U9645 ( .A(n9838), .B(n9839), .Z(n9640) );
  ANDN U9646 ( .A(n9840), .B(n9841), .Z(n9839) );
  XNOR U9647 ( .A(n9838), .B(n9842), .Z(n9840) );
  XOR U9648 ( .A(n9650), .B(n9843), .Z(n9644) );
  IV U9649 ( .A(n9649), .Z(n9843) );
  XNOR U9650 ( .A(n9646), .B(n9798), .Z(n9649) );
  AND U9651 ( .A(n11049), .B(n8272), .Z(n9798) );
  XOR U9652 ( .A(n9844), .B(n9845), .Z(n9646) );
  ANDN U9653 ( .A(n9846), .B(n9847), .Z(n9845) );
  XNOR U9654 ( .A(n9844), .B(n9848), .Z(n9846) );
  XOR U9655 ( .A(n9656), .B(n9849), .Z(n9650) );
  IV U9656 ( .A(n9655), .Z(n9849) );
  XNOR U9657 ( .A(n9652), .B(n9791), .Z(n9655) );
  AND U9658 ( .A(n11341), .B(n7770), .Z(n9791) );
  XOR U9659 ( .A(n9850), .B(n9851), .Z(n9652) );
  ANDN U9660 ( .A(n9852), .B(n9853), .Z(n9851) );
  XNOR U9661 ( .A(n9850), .B(n9854), .Z(n9852) );
  XOR U9662 ( .A(n9662), .B(n9855), .Z(n9656) );
  IV U9663 ( .A(n9661), .Z(n9855) );
  XNOR U9664 ( .A(n9658), .B(n9784), .Z(n9661) );
  AND U9665 ( .A(n11607), .B(n7241), .Z(n9784) );
  XOR U9666 ( .A(n9856), .B(n9857), .Z(n9658) );
  ANDN U9667 ( .A(n9858), .B(n9859), .Z(n9857) );
  XNOR U9668 ( .A(n9856), .B(n9860), .Z(n9858) );
  XOR U9669 ( .A(n9668), .B(n9861), .Z(n9662) );
  IV U9670 ( .A(n9667), .Z(n9861) );
  XNOR U9671 ( .A(n9664), .B(n9777), .Z(n9667) );
  AND U9672 ( .A(n11869), .B(n6688), .Z(n9777) );
  XOR U9673 ( .A(n9862), .B(n9863), .Z(n9664) );
  ANDN U9674 ( .A(n9864), .B(n9865), .Z(n9863) );
  XNOR U9675 ( .A(n9862), .B(n9866), .Z(n9864) );
  XOR U9676 ( .A(n9674), .B(n9867), .Z(n9668) );
  IV U9677 ( .A(n9673), .Z(n9867) );
  XNOR U9678 ( .A(n9670), .B(n9770), .Z(n9673) );
  AND U9679 ( .A(n12128), .B(n6118), .Z(n9770) );
  XOR U9680 ( .A(n9868), .B(n9869), .Z(n9670) );
  ANDN U9681 ( .A(n9870), .B(n9871), .Z(n9869) );
  XNOR U9682 ( .A(n9868), .B(n9872), .Z(n9870) );
  XOR U9683 ( .A(n9680), .B(n9873), .Z(n9674) );
  IV U9684 ( .A(n9679), .Z(n9873) );
  XNOR U9685 ( .A(n9676), .B(n9763), .Z(n9679) );
  AND U9686 ( .A(n12387), .B(n5561), .Z(n9763) );
  XOR U9687 ( .A(n9874), .B(n9875), .Z(n9676) );
  ANDN U9688 ( .A(n9876), .B(n9877), .Z(n9875) );
  XNOR U9689 ( .A(n9874), .B(n9878), .Z(n9876) );
  XOR U9690 ( .A(n9686), .B(n9879), .Z(n9680) );
  IV U9691 ( .A(n9685), .Z(n9879) );
  XNOR U9692 ( .A(n9682), .B(n9756), .Z(n9685) );
  AND U9693 ( .A(n12644), .B(n5030), .Z(n9756) );
  XOR U9694 ( .A(n9880), .B(n9881), .Z(n9682) );
  ANDN U9695 ( .A(n9882), .B(n9883), .Z(n9881) );
  XNOR U9696 ( .A(n9880), .B(n9884), .Z(n9882) );
  XOR U9697 ( .A(n9692), .B(n9885), .Z(n9686) );
  IV U9698 ( .A(n9691), .Z(n9885) );
  XNOR U9699 ( .A(n9688), .B(n9749), .Z(n9691) );
  AND U9700 ( .A(n12880), .B(n4525), .Z(n9749) );
  XOR U9701 ( .A(n9886), .B(n9887), .Z(n9688) );
  ANDN U9702 ( .A(n9888), .B(n9889), .Z(n9887) );
  XNOR U9703 ( .A(n9886), .B(n9890), .Z(n9888) );
  XOR U9704 ( .A(n9698), .B(n9891), .Z(n9692) );
  IV U9705 ( .A(n9697), .Z(n9891) );
  XNOR U9706 ( .A(n9694), .B(n9742), .Z(n9697) );
  AND U9707 ( .A(n13070), .B(n4046), .Z(n9742) );
  XOR U9708 ( .A(n9892), .B(n9893), .Z(n9694) );
  ANDN U9709 ( .A(n9894), .B(n9895), .Z(n9893) );
  XNOR U9710 ( .A(n9892), .B(n9896), .Z(n9894) );
  XOR U9711 ( .A(n9704), .B(n9897), .Z(n9698) );
  IV U9712 ( .A(n9703), .Z(n9897) );
  XNOR U9713 ( .A(n9700), .B(n9735), .Z(n9703) );
  AND U9714 ( .A(n13207), .B(n3593), .Z(n9735) );
  XOR U9715 ( .A(n9898), .B(n9899), .Z(n9700) );
  ANDN U9716 ( .A(n9900), .B(n9901), .Z(n9899) );
  XNOR U9717 ( .A(n9898), .B(n9902), .Z(n9900) );
  XNOR U9718 ( .A(n9709), .B(n9527), .Z(n9704) );
  XNOR U9719 ( .A(n9706), .B(n9903), .Z(n9709) );
  AND U9720 ( .A(n6527), .B(n3166), .Z(n9903) );
  XOR U9721 ( .A(n9904), .B(n9905), .Z(n9706) );
  ANDN U9722 ( .A(n9906), .B(n9907), .Z(n9905) );
  XNOR U9723 ( .A(n9732), .B(n9904), .Z(n9906) );
  XOR U9724 ( .A(n9908), .B(n9527), .Z(n9729) );
  NANDN U9725 ( .B(n6808), .A(n2765), .Z(n9527) );
  XOR U9726 ( .A(n9909), .B(n9910), .Z(n2765) );
  AND U9727 ( .A(n6809), .B(n9911), .Z(n9910) );
  XNOR U9728 ( .A(n9909), .B(n9716), .Z(n9911) );
  XOR U9729 ( .A(n9714), .B(n9909), .Z(n9716) );
  XOR U9730 ( .A(n9912), .B(n9913), .Z(n9714) );
  ANDN U9731 ( .A(n9912), .B(n9914), .Z(n9913) );
  XOR U9732 ( .A(n9915), .B(n7368), .Z(n9909) );
  IV U9733 ( .A(n9718), .Z(n9908) );
  XOR U9734 ( .A(n9916), .B(n9917), .Z(n9718) );
  AND U9735 ( .A(n9918), .B(n9919), .Z(n9917) );
  XNOR U9736 ( .A(n9920), .B(n9916), .Z(n9919) );
  XNOR U9737 ( .A(n9722), .B(n9725), .Z(n9728) );
  XOR U9738 ( .A(n9921), .B(n9922), .Z(n9722) );
  XOR U9739 ( .A(n9923), .B(n9924), .Z(n9725) );
  AND U9740 ( .A(n9923), .B(n9925), .Z(n9924) );
  XOR U9741 ( .A(n9926), .B(n9918), .Z(n9925) );
  XOR U9742 ( .A(n9927), .B(n9733), .Z(n9918) );
  XOR U9743 ( .A(n9740), .B(n9928), .Z(n9733) );
  IV U9744 ( .A(n9738), .Z(n9928) );
  XNOR U9745 ( .A(n9929), .B(n9737), .Z(n9738) );
  OR U9746 ( .A(n9930), .B(n9931), .Z(n9737) );
  NANDN U9747 ( .B(n6541), .A(n3593), .Z(n9929) );
  XOR U9748 ( .A(n9747), .B(n9932), .Z(n9740) );
  IV U9749 ( .A(n9746), .Z(n9932) );
  XNOR U9750 ( .A(n9743), .B(n9933), .Z(n9746) );
  XOR U9751 ( .A(n9934), .B(n9935), .Z(n9743) );
  NANDN U9752 ( .B(n9936), .A(n9937), .Z(n9934) );
  XOR U9753 ( .A(n9935), .B(n9938), .Z(n9937) );
  XOR U9754 ( .A(n9754), .B(n9939), .Z(n9747) );
  IV U9755 ( .A(n9753), .Z(n9939) );
  XNOR U9756 ( .A(n9750), .B(n9940), .Z(n9753) );
  XOR U9757 ( .A(n9941), .B(n9942), .Z(n9750) );
  ANDN U9758 ( .A(n9943), .B(n9944), .Z(n9942) );
  XNOR U9759 ( .A(n9941), .B(n9945), .Z(n9943) );
  XOR U9760 ( .A(n9761), .B(n9946), .Z(n9754) );
  IV U9761 ( .A(n9760), .Z(n9946) );
  XNOR U9762 ( .A(n9757), .B(n9947), .Z(n9760) );
  XOR U9763 ( .A(n9948), .B(n9949), .Z(n9757) );
  ANDN U9764 ( .A(n9950), .B(n9951), .Z(n9949) );
  XNOR U9765 ( .A(n9948), .B(n9952), .Z(n9950) );
  XOR U9766 ( .A(n9768), .B(n9953), .Z(n9761) );
  IV U9767 ( .A(n9767), .Z(n9953) );
  XNOR U9768 ( .A(n9764), .B(n9954), .Z(n9767) );
  XOR U9769 ( .A(n9955), .B(n9956), .Z(n9764) );
  ANDN U9770 ( .A(n9957), .B(n9958), .Z(n9956) );
  XNOR U9771 ( .A(n9955), .B(n9959), .Z(n9957) );
  XOR U9772 ( .A(n9775), .B(n9960), .Z(n9768) );
  IV U9773 ( .A(n9774), .Z(n9960) );
  XNOR U9774 ( .A(n9771), .B(n9961), .Z(n9774) );
  XOR U9775 ( .A(n9962), .B(n9963), .Z(n9771) );
  ANDN U9776 ( .A(n9964), .B(n9965), .Z(n9963) );
  XNOR U9777 ( .A(n9962), .B(n9966), .Z(n9964) );
  XOR U9778 ( .A(n9782), .B(n9967), .Z(n9775) );
  IV U9779 ( .A(n9781), .Z(n9967) );
  XNOR U9780 ( .A(n9778), .B(n9968), .Z(n9781) );
  XOR U9781 ( .A(n9969), .B(n9970), .Z(n9778) );
  ANDN U9782 ( .A(n9971), .B(n9972), .Z(n9970) );
  XNOR U9783 ( .A(n9969), .B(n9973), .Z(n9971) );
  XOR U9784 ( .A(n9789), .B(n9974), .Z(n9782) );
  IV U9785 ( .A(n9788), .Z(n9974) );
  XNOR U9786 ( .A(n9785), .B(n9975), .Z(n9788) );
  XOR U9787 ( .A(n9976), .B(n9977), .Z(n9785) );
  ANDN U9788 ( .A(n9978), .B(n9979), .Z(n9977) );
  XNOR U9789 ( .A(n9976), .B(n9980), .Z(n9978) );
  XOR U9790 ( .A(n9796), .B(n9981), .Z(n9789) );
  IV U9791 ( .A(n9795), .Z(n9981) );
  XNOR U9792 ( .A(n9792), .B(n9982), .Z(n9795) );
  XOR U9793 ( .A(n9983), .B(n9984), .Z(n9792) );
  ANDN U9794 ( .A(n9985), .B(n9986), .Z(n9984) );
  XNOR U9795 ( .A(n9983), .B(n9987), .Z(n9985) );
  XOR U9796 ( .A(n9803), .B(n9988), .Z(n9796) );
  IV U9797 ( .A(n9802), .Z(n9988) );
  XNOR U9798 ( .A(n9799), .B(n9989), .Z(n9802) );
  XOR U9799 ( .A(n9990), .B(n9991), .Z(n9799) );
  ANDN U9800 ( .A(n9992), .B(n9993), .Z(n9991) );
  XNOR U9801 ( .A(n9990), .B(n9994), .Z(n9992) );
  XOR U9802 ( .A(n9810), .B(n9995), .Z(n9803) );
  IV U9803 ( .A(n9809), .Z(n9995) );
  XNOR U9804 ( .A(n9806), .B(n9996), .Z(n9809) );
  XOR U9805 ( .A(n9997), .B(n9998), .Z(n9806) );
  ANDN U9806 ( .A(n9999), .B(n10000), .Z(n9998) );
  XNOR U9807 ( .A(n9997), .B(n10001), .Z(n9999) );
  XOR U9808 ( .A(n9817), .B(n10002), .Z(n9810) );
  IV U9809 ( .A(n9816), .Z(n10002) );
  XNOR U9810 ( .A(n9813), .B(n10003), .Z(n9816) );
  XOR U9811 ( .A(n10004), .B(n10005), .Z(n9813) );
  ANDN U9812 ( .A(n10006), .B(n10007), .Z(n10005) );
  XNOR U9813 ( .A(n10004), .B(n10008), .Z(n10006) );
  XOR U9814 ( .A(n9824), .B(n10009), .Z(n9817) );
  IV U9815 ( .A(n9823), .Z(n10009) );
  XNOR U9816 ( .A(n9820), .B(n10010), .Z(n9823) );
  XOR U9817 ( .A(n10011), .B(n10012), .Z(n9820) );
  ANDN U9818 ( .A(n10013), .B(n10014), .Z(n10012) );
  XNOR U9819 ( .A(n10011), .B(n10015), .Z(n10013) );
  XOR U9820 ( .A(n9830), .B(n10016), .Z(n9824) );
  IV U9821 ( .A(n9829), .Z(n10016) );
  XNOR U9822 ( .A(n9826), .B(n10017), .Z(n9829) );
  XOR U9823 ( .A(n10018), .B(n10019), .Z(n9826) );
  ANDN U9824 ( .A(n10020), .B(n10021), .Z(n10019) );
  XNOR U9825 ( .A(n10018), .B(n10022), .Z(n10020) );
  XOR U9826 ( .A(n9836), .B(n10023), .Z(n9830) );
  IV U9827 ( .A(n9835), .Z(n10023) );
  XNOR U9828 ( .A(n9832), .B(n10010), .Z(n9835) );
  AND U9829 ( .A(n10387), .B(n9621), .Z(n10010) );
  XOR U9830 ( .A(n10024), .B(n10025), .Z(n9832) );
  ANDN U9831 ( .A(n10026), .B(n10027), .Z(n10025) );
  XNOR U9832 ( .A(n10024), .B(n10028), .Z(n10026) );
  XOR U9833 ( .A(n9842), .B(n10029), .Z(n9836) );
  IV U9834 ( .A(n9841), .Z(n10029) );
  XNOR U9835 ( .A(n9838), .B(n10003), .Z(n9841) );
  AND U9836 ( .A(n10731), .B(n9198), .Z(n10003) );
  XOR U9837 ( .A(n10030), .B(n10031), .Z(n9838) );
  ANDN U9838 ( .A(n10032), .B(n10033), .Z(n10031) );
  XNOR U9839 ( .A(n10030), .B(n10034), .Z(n10032) );
  XOR U9840 ( .A(n9848), .B(n10035), .Z(n9842) );
  IV U9841 ( .A(n9847), .Z(n10035) );
  XNOR U9842 ( .A(n9844), .B(n9996), .Z(n9847) );
  AND U9843 ( .A(n11049), .B(n8748), .Z(n9996) );
  XOR U9844 ( .A(n10036), .B(n10037), .Z(n9844) );
  ANDN U9845 ( .A(n10038), .B(n10039), .Z(n10037) );
  XNOR U9846 ( .A(n10036), .B(n10040), .Z(n10038) );
  XOR U9847 ( .A(n9854), .B(n10041), .Z(n9848) );
  IV U9848 ( .A(n9853), .Z(n10041) );
  XNOR U9849 ( .A(n9850), .B(n9989), .Z(n9853) );
  AND U9850 ( .A(n11341), .B(n8272), .Z(n9989) );
  XOR U9851 ( .A(n10042), .B(n10043), .Z(n9850) );
  ANDN U9852 ( .A(n10044), .B(n10045), .Z(n10043) );
  XNOR U9853 ( .A(n10042), .B(n10046), .Z(n10044) );
  XOR U9854 ( .A(n9860), .B(n10047), .Z(n9854) );
  IV U9855 ( .A(n9859), .Z(n10047) );
  XNOR U9856 ( .A(n9856), .B(n9982), .Z(n9859) );
  AND U9857 ( .A(n11607), .B(n7770), .Z(n9982) );
  XOR U9858 ( .A(n10048), .B(n10049), .Z(n9856) );
  ANDN U9859 ( .A(n10050), .B(n10051), .Z(n10049) );
  XNOR U9860 ( .A(n10048), .B(n10052), .Z(n10050) );
  XOR U9861 ( .A(n9866), .B(n10053), .Z(n9860) );
  IV U9862 ( .A(n9865), .Z(n10053) );
  XNOR U9863 ( .A(n9862), .B(n9975), .Z(n9865) );
  AND U9864 ( .A(n11869), .B(n7241), .Z(n9975) );
  XOR U9865 ( .A(n10054), .B(n10055), .Z(n9862) );
  ANDN U9866 ( .A(n10056), .B(n10057), .Z(n10055) );
  XNOR U9867 ( .A(n10054), .B(n10058), .Z(n10056) );
  XOR U9868 ( .A(n9872), .B(n10059), .Z(n9866) );
  IV U9869 ( .A(n9871), .Z(n10059) );
  XNOR U9870 ( .A(n9868), .B(n9968), .Z(n9871) );
  AND U9871 ( .A(n12128), .B(n6688), .Z(n9968) );
  XOR U9872 ( .A(n10060), .B(n10061), .Z(n9868) );
  ANDN U9873 ( .A(n10062), .B(n10063), .Z(n10061) );
  XNOR U9874 ( .A(n10060), .B(n10064), .Z(n10062) );
  XOR U9875 ( .A(n9878), .B(n10065), .Z(n9872) );
  IV U9876 ( .A(n9877), .Z(n10065) );
  XNOR U9877 ( .A(n9874), .B(n9961), .Z(n9877) );
  AND U9878 ( .A(n12387), .B(n6118), .Z(n9961) );
  XOR U9879 ( .A(n10066), .B(n10067), .Z(n9874) );
  ANDN U9880 ( .A(n10068), .B(n10069), .Z(n10067) );
  XNOR U9881 ( .A(n10066), .B(n10070), .Z(n10068) );
  XOR U9882 ( .A(n9884), .B(n10071), .Z(n9878) );
  IV U9883 ( .A(n9883), .Z(n10071) );
  XNOR U9884 ( .A(n9880), .B(n9954), .Z(n9883) );
  AND U9885 ( .A(n12644), .B(n5561), .Z(n9954) );
  XOR U9886 ( .A(n10072), .B(n10073), .Z(n9880) );
  ANDN U9887 ( .A(n10074), .B(n10075), .Z(n10073) );
  XNOR U9888 ( .A(n10072), .B(n10076), .Z(n10074) );
  XOR U9889 ( .A(n9890), .B(n10077), .Z(n9884) );
  IV U9890 ( .A(n9889), .Z(n10077) );
  XNOR U9891 ( .A(n9886), .B(n9947), .Z(n9889) );
  AND U9892 ( .A(n12880), .B(n5030), .Z(n9947) );
  XOR U9893 ( .A(n10078), .B(n10079), .Z(n9886) );
  ANDN U9894 ( .A(n10080), .B(n10081), .Z(n10079) );
  XNOR U9895 ( .A(n10078), .B(n10082), .Z(n10080) );
  XOR U9896 ( .A(n9896), .B(n10083), .Z(n9890) );
  IV U9897 ( .A(n9895), .Z(n10083) );
  XNOR U9898 ( .A(n9892), .B(n9940), .Z(n9895) );
  AND U9899 ( .A(n13070), .B(n4525), .Z(n9940) );
  XOR U9900 ( .A(n10084), .B(n10085), .Z(n9892) );
  ANDN U9901 ( .A(n10086), .B(n10087), .Z(n10085) );
  XNOR U9902 ( .A(n10084), .B(n10088), .Z(n10086) );
  XOR U9903 ( .A(n9902), .B(n10089), .Z(n9896) );
  IV U9904 ( .A(n9901), .Z(n10089) );
  XNOR U9905 ( .A(n9898), .B(n9933), .Z(n9901) );
  AND U9906 ( .A(n13207), .B(n4046), .Z(n9933) );
  XOR U9907 ( .A(n10090), .B(n10091), .Z(n9898) );
  ANDN U9908 ( .A(n10092), .B(n10093), .Z(n10091) );
  XNOR U9909 ( .A(n10090), .B(n10094), .Z(n10092) );
  XNOR U9910 ( .A(n9907), .B(n9732), .Z(n9902) );
  XNOR U9911 ( .A(n9904), .B(n10095), .Z(n9907) );
  AND U9912 ( .A(n6527), .B(n3593), .Z(n10095) );
  XOR U9913 ( .A(n10096), .B(n10097), .Z(n9904) );
  ANDN U9914 ( .A(n10098), .B(n10099), .Z(n10097) );
  XNOR U9915 ( .A(n9930), .B(n10096), .Z(n10098) );
  XOR U9916 ( .A(n10100), .B(n9732), .Z(n9927) );
  NANDN U9917 ( .B(n6808), .A(n3166), .Z(n9732) );
  XOR U9918 ( .A(n10101), .B(n10102), .Z(n3166) );
  AND U9919 ( .A(n6809), .B(n10103), .Z(n10102) );
  XNOR U9920 ( .A(n10101), .B(n9914), .Z(n10103) );
  XOR U9921 ( .A(n9912), .B(n10101), .Z(n9914) );
  XOR U9922 ( .A(n10104), .B(n10105), .Z(n9912) );
  ANDN U9923 ( .A(n10104), .B(n10106), .Z(n10105) );
  XOR U9924 ( .A(n10107), .B(n7368), .Z(n10101) );
  IV U9925 ( .A(n9916), .Z(n10100) );
  XOR U9926 ( .A(n10108), .B(n10109), .Z(n9916) );
  AND U9927 ( .A(n10110), .B(n10111), .Z(n10109) );
  XNOR U9928 ( .A(n10112), .B(n10108), .Z(n10111) );
  XNOR U9929 ( .A(n9920), .B(n9923), .Z(n9926) );
  XOR U9930 ( .A(n10113), .B(n10114), .Z(n9920) );
  XOR U9931 ( .A(n10115), .B(n10116), .Z(n9923) );
  AND U9932 ( .A(n10115), .B(n10117), .Z(n10116) );
  XOR U9933 ( .A(n10118), .B(n10110), .Z(n10117) );
  XOR U9934 ( .A(n10119), .B(n9931), .Z(n10110) );
  XOR U9935 ( .A(n9938), .B(n10120), .Z(n9931) );
  IV U9936 ( .A(n9936), .Z(n10120) );
  XNOR U9937 ( .A(n10121), .B(n9935), .Z(n9936) );
  OR U9938 ( .A(n10122), .B(n10123), .Z(n9935) );
  NANDN U9939 ( .B(n6541), .A(n4046), .Z(n10121) );
  XOR U9940 ( .A(n9945), .B(n10124), .Z(n9938) );
  IV U9941 ( .A(n9944), .Z(n10124) );
  XNOR U9942 ( .A(n9941), .B(n10125), .Z(n9944) );
  XOR U9943 ( .A(n10126), .B(n10127), .Z(n9941) );
  NANDN U9944 ( .B(n10128), .A(n10129), .Z(n10126) );
  XOR U9945 ( .A(n10127), .B(n10130), .Z(n10129) );
  XOR U9946 ( .A(n9952), .B(n10131), .Z(n9945) );
  IV U9947 ( .A(n9951), .Z(n10131) );
  XNOR U9948 ( .A(n9948), .B(n10132), .Z(n9951) );
  XOR U9949 ( .A(n10133), .B(n10134), .Z(n9948) );
  ANDN U9950 ( .A(n10135), .B(n10136), .Z(n10134) );
  XNOR U9951 ( .A(n10133), .B(n10137), .Z(n10135) );
  XOR U9952 ( .A(n9959), .B(n10138), .Z(n9952) );
  IV U9953 ( .A(n9958), .Z(n10138) );
  XNOR U9954 ( .A(n9955), .B(n10139), .Z(n9958) );
  XOR U9955 ( .A(n10140), .B(n10141), .Z(n9955) );
  ANDN U9956 ( .A(n10142), .B(n10143), .Z(n10141) );
  XNOR U9957 ( .A(n10140), .B(n10144), .Z(n10142) );
  XOR U9958 ( .A(n9966), .B(n10145), .Z(n9959) );
  IV U9959 ( .A(n9965), .Z(n10145) );
  XNOR U9960 ( .A(n9962), .B(n10146), .Z(n9965) );
  XOR U9961 ( .A(n10147), .B(n10148), .Z(n9962) );
  ANDN U9962 ( .A(n10149), .B(n10150), .Z(n10148) );
  XNOR U9963 ( .A(n10147), .B(n10151), .Z(n10149) );
  XOR U9964 ( .A(n9973), .B(n10152), .Z(n9966) );
  IV U9965 ( .A(n9972), .Z(n10152) );
  XNOR U9966 ( .A(n9969), .B(n10153), .Z(n9972) );
  XOR U9967 ( .A(n10154), .B(n10155), .Z(n9969) );
  ANDN U9968 ( .A(n10156), .B(n10157), .Z(n10155) );
  XNOR U9969 ( .A(n10154), .B(n10158), .Z(n10156) );
  XOR U9970 ( .A(n9980), .B(n10159), .Z(n9973) );
  IV U9971 ( .A(n9979), .Z(n10159) );
  XNOR U9972 ( .A(n9976), .B(n10160), .Z(n9979) );
  XOR U9973 ( .A(n10161), .B(n10162), .Z(n9976) );
  ANDN U9974 ( .A(n10163), .B(n10164), .Z(n10162) );
  XNOR U9975 ( .A(n10161), .B(n10165), .Z(n10163) );
  XOR U9976 ( .A(n9987), .B(n10166), .Z(n9980) );
  IV U9977 ( .A(n9986), .Z(n10166) );
  XNOR U9978 ( .A(n9983), .B(n10167), .Z(n9986) );
  XOR U9979 ( .A(n10168), .B(n10169), .Z(n9983) );
  ANDN U9980 ( .A(n10170), .B(n10171), .Z(n10169) );
  XNOR U9981 ( .A(n10168), .B(n10172), .Z(n10170) );
  XOR U9982 ( .A(n9994), .B(n10173), .Z(n9987) );
  IV U9983 ( .A(n9993), .Z(n10173) );
  XNOR U9984 ( .A(n9990), .B(n10174), .Z(n9993) );
  XOR U9985 ( .A(n10175), .B(n10176), .Z(n9990) );
  ANDN U9986 ( .A(n10177), .B(n10178), .Z(n10176) );
  XNOR U9987 ( .A(n10175), .B(n10179), .Z(n10177) );
  XOR U9988 ( .A(n10001), .B(n10180), .Z(n9994) );
  IV U9989 ( .A(n10000), .Z(n10180) );
  XNOR U9990 ( .A(n9997), .B(n10181), .Z(n10000) );
  XOR U9991 ( .A(n10182), .B(n10183), .Z(n9997) );
  ANDN U9992 ( .A(n10184), .B(n10185), .Z(n10183) );
  XNOR U9993 ( .A(n10182), .B(n10186), .Z(n10184) );
  XOR U9994 ( .A(n10008), .B(n10187), .Z(n10001) );
  IV U9995 ( .A(n10007), .Z(n10187) );
  XNOR U9996 ( .A(n10004), .B(n10188), .Z(n10007) );
  XOR U9997 ( .A(n10189), .B(n10190), .Z(n10004) );
  ANDN U9998 ( .A(n10191), .B(n10192), .Z(n10190) );
  XNOR U9999 ( .A(n10189), .B(n10193), .Z(n10191) );
  XOR U10000 ( .A(n10015), .B(n10194), .Z(n10008) );
  IV U10001 ( .A(n10014), .Z(n10194) );
  XNOR U10002 ( .A(n10011), .B(n10195), .Z(n10014) );
  XOR U10003 ( .A(n10196), .B(n10197), .Z(n10011) );
  ANDN U10004 ( .A(n10198), .B(n10199), .Z(n10197) );
  XNOR U10005 ( .A(n10196), .B(n10200), .Z(n10198) );
  XOR U10006 ( .A(n10022), .B(n10201), .Z(n10015) );
  IV U10007 ( .A(n10021), .Z(n10201) );
  XNOR U10008 ( .A(n10018), .B(n10202), .Z(n10021) );
  XOR U10009 ( .A(n10203), .B(n10204), .Z(n10018) );
  ANDN U10010 ( .A(n10205), .B(n10206), .Z(n10204) );
  XNOR U10011 ( .A(n10203), .B(n10207), .Z(n10205) );
  XOR U10012 ( .A(n10028), .B(n10208), .Z(n10022) );
  IV U10013 ( .A(n10027), .Z(n10208) );
  XNOR U10014 ( .A(n10024), .B(n10202), .Z(n10027) );
  AND U10015 ( .A(n10387), .B(n10017), .Z(n10202) );
  XOR U10016 ( .A(n10209), .B(n10210), .Z(n10024) );
  ANDN U10017 ( .A(n10211), .B(n10212), .Z(n10210) );
  XNOR U10018 ( .A(n10209), .B(n10213), .Z(n10211) );
  XOR U10019 ( .A(n10034), .B(n10214), .Z(n10028) );
  IV U10020 ( .A(n10033), .Z(n10214) );
  XNOR U10021 ( .A(n10030), .B(n10195), .Z(n10033) );
  AND U10022 ( .A(n10731), .B(n9621), .Z(n10195) );
  XOR U10023 ( .A(n10215), .B(n10216), .Z(n10030) );
  ANDN U10024 ( .A(n10217), .B(n10218), .Z(n10216) );
  XNOR U10025 ( .A(n10215), .B(n10219), .Z(n10217) );
  XOR U10026 ( .A(n10040), .B(n10220), .Z(n10034) );
  IV U10027 ( .A(n10039), .Z(n10220) );
  XNOR U10028 ( .A(n10036), .B(n10188), .Z(n10039) );
  AND U10029 ( .A(n11049), .B(n9198), .Z(n10188) );
  XOR U10030 ( .A(n10221), .B(n10222), .Z(n10036) );
  ANDN U10031 ( .A(n10223), .B(n10224), .Z(n10222) );
  XNOR U10032 ( .A(n10221), .B(n10225), .Z(n10223) );
  XOR U10033 ( .A(n10046), .B(n10226), .Z(n10040) );
  IV U10034 ( .A(n10045), .Z(n10226) );
  XNOR U10035 ( .A(n10042), .B(n10181), .Z(n10045) );
  AND U10036 ( .A(n11341), .B(n8748), .Z(n10181) );
  XOR U10037 ( .A(n10227), .B(n10228), .Z(n10042) );
  ANDN U10038 ( .A(n10229), .B(n10230), .Z(n10228) );
  XNOR U10039 ( .A(n10227), .B(n10231), .Z(n10229) );
  XOR U10040 ( .A(n10052), .B(n10232), .Z(n10046) );
  IV U10041 ( .A(n10051), .Z(n10232) );
  XNOR U10042 ( .A(n10048), .B(n10174), .Z(n10051) );
  AND U10043 ( .A(n11607), .B(n8272), .Z(n10174) );
  XOR U10044 ( .A(n10233), .B(n10234), .Z(n10048) );
  ANDN U10045 ( .A(n10235), .B(n10236), .Z(n10234) );
  XNOR U10046 ( .A(n10233), .B(n10237), .Z(n10235) );
  XOR U10047 ( .A(n10058), .B(n10238), .Z(n10052) );
  IV U10048 ( .A(n10057), .Z(n10238) );
  XNOR U10049 ( .A(n10054), .B(n10167), .Z(n10057) );
  AND U10050 ( .A(n11869), .B(n7770), .Z(n10167) );
  XOR U10051 ( .A(n10239), .B(n10240), .Z(n10054) );
  ANDN U10052 ( .A(n10241), .B(n10242), .Z(n10240) );
  XNOR U10053 ( .A(n10239), .B(n10243), .Z(n10241) );
  XOR U10054 ( .A(n10064), .B(n10244), .Z(n10058) );
  IV U10055 ( .A(n10063), .Z(n10244) );
  XNOR U10056 ( .A(n10060), .B(n10160), .Z(n10063) );
  AND U10057 ( .A(n12128), .B(n7241), .Z(n10160) );
  XOR U10058 ( .A(n10245), .B(n10246), .Z(n10060) );
  ANDN U10059 ( .A(n10247), .B(n10248), .Z(n10246) );
  XNOR U10060 ( .A(n10245), .B(n10249), .Z(n10247) );
  XOR U10061 ( .A(n10070), .B(n10250), .Z(n10064) );
  IV U10062 ( .A(n10069), .Z(n10250) );
  XNOR U10063 ( .A(n10066), .B(n10153), .Z(n10069) );
  AND U10064 ( .A(n12387), .B(n6688), .Z(n10153) );
  XOR U10065 ( .A(n10251), .B(n10252), .Z(n10066) );
  ANDN U10066 ( .A(n10253), .B(n10254), .Z(n10252) );
  XNOR U10067 ( .A(n10251), .B(n10255), .Z(n10253) );
  XOR U10068 ( .A(n10076), .B(n10256), .Z(n10070) );
  IV U10069 ( .A(n10075), .Z(n10256) );
  XNOR U10070 ( .A(n10072), .B(n10146), .Z(n10075) );
  AND U10071 ( .A(n12644), .B(n6118), .Z(n10146) );
  XOR U10072 ( .A(n10257), .B(n10258), .Z(n10072) );
  ANDN U10073 ( .A(n10259), .B(n10260), .Z(n10258) );
  XNOR U10074 ( .A(n10257), .B(n10261), .Z(n10259) );
  XOR U10075 ( .A(n10082), .B(n10262), .Z(n10076) );
  IV U10076 ( .A(n10081), .Z(n10262) );
  XNOR U10077 ( .A(n10078), .B(n10139), .Z(n10081) );
  AND U10078 ( .A(n12880), .B(n5561), .Z(n10139) );
  XOR U10079 ( .A(n10263), .B(n10264), .Z(n10078) );
  ANDN U10080 ( .A(n10265), .B(n10266), .Z(n10264) );
  XNOR U10081 ( .A(n10263), .B(n10267), .Z(n10265) );
  XOR U10082 ( .A(n10088), .B(n10268), .Z(n10082) );
  IV U10083 ( .A(n10087), .Z(n10268) );
  XNOR U10084 ( .A(n10084), .B(n10132), .Z(n10087) );
  AND U10085 ( .A(n13070), .B(n5030), .Z(n10132) );
  XOR U10086 ( .A(n10269), .B(n10270), .Z(n10084) );
  ANDN U10087 ( .A(n10271), .B(n10272), .Z(n10270) );
  XNOR U10088 ( .A(n10269), .B(n10273), .Z(n10271) );
  XOR U10089 ( .A(n10094), .B(n10274), .Z(n10088) );
  IV U10090 ( .A(n10093), .Z(n10274) );
  XNOR U10091 ( .A(n10090), .B(n10125), .Z(n10093) );
  AND U10092 ( .A(n13207), .B(n4525), .Z(n10125) );
  XOR U10093 ( .A(n10275), .B(n10276), .Z(n10090) );
  ANDN U10094 ( .A(n10277), .B(n10278), .Z(n10276) );
  XNOR U10095 ( .A(n10275), .B(n10279), .Z(n10277) );
  XNOR U10096 ( .A(n10099), .B(n9930), .Z(n10094) );
  XNOR U10097 ( .A(n10096), .B(n10280), .Z(n10099) );
  AND U10098 ( .A(n6527), .B(n4046), .Z(n10280) );
  XOR U10099 ( .A(n10281), .B(n10282), .Z(n10096) );
  ANDN U10100 ( .A(n10283), .B(n10284), .Z(n10282) );
  XNOR U10101 ( .A(n10122), .B(n10281), .Z(n10283) );
  XOR U10102 ( .A(n10285), .B(n9930), .Z(n10119) );
  NANDN U10103 ( .B(n6808), .A(n3593), .Z(n9930) );
  XOR U10104 ( .A(n10286), .B(n10287), .Z(n3593) );
  AND U10105 ( .A(n6809), .B(n10288), .Z(n10287) );
  XNOR U10106 ( .A(n10286), .B(n10106), .Z(n10288) );
  XOR U10107 ( .A(n10104), .B(n10286), .Z(n10106) );
  XOR U10108 ( .A(n10289), .B(n10290), .Z(n10104) );
  ANDN U10109 ( .A(n10289), .B(n10291), .Z(n10290) );
  XOR U10110 ( .A(n10292), .B(n7368), .Z(n10286) );
  IV U10111 ( .A(n10108), .Z(n10285) );
  XOR U10112 ( .A(n10293), .B(n10294), .Z(n10108) );
  AND U10113 ( .A(n10295), .B(n10296), .Z(n10294) );
  XNOR U10114 ( .A(n10297), .B(n10293), .Z(n10296) );
  XNOR U10115 ( .A(n10112), .B(n10115), .Z(n10118) );
  XOR U10116 ( .A(n10298), .B(n10299), .Z(n10112) );
  XOR U10117 ( .A(n10300), .B(n10301), .Z(n10115) );
  AND U10118 ( .A(n10300), .B(n10302), .Z(n10301) );
  XOR U10119 ( .A(n10303), .B(n10295), .Z(n10302) );
  XOR U10120 ( .A(n10304), .B(n10123), .Z(n10295) );
  XOR U10121 ( .A(n10130), .B(n10305), .Z(n10123) );
  IV U10122 ( .A(n10128), .Z(n10305) );
  XNOR U10123 ( .A(n10306), .B(n10127), .Z(n10128) );
  OR U10124 ( .A(n10307), .B(n10308), .Z(n10127) );
  NANDN U10125 ( .B(n6541), .A(n4525), .Z(n10306) );
  XOR U10126 ( .A(n10137), .B(n10309), .Z(n10130) );
  IV U10127 ( .A(n10136), .Z(n10309) );
  XNOR U10128 ( .A(n10133), .B(n10310), .Z(n10136) );
  XOR U10129 ( .A(n10311), .B(n10312), .Z(n10133) );
  NANDN U10130 ( .B(n10313), .A(n10314), .Z(n10311) );
  XOR U10131 ( .A(n10312), .B(n10315), .Z(n10314) );
  XOR U10132 ( .A(n10144), .B(n10316), .Z(n10137) );
  IV U10133 ( .A(n10143), .Z(n10316) );
  XNOR U10134 ( .A(n10140), .B(n10317), .Z(n10143) );
  XOR U10135 ( .A(n10318), .B(n10319), .Z(n10140) );
  ANDN U10136 ( .A(n10320), .B(n10321), .Z(n10319) );
  XNOR U10137 ( .A(n10318), .B(n10322), .Z(n10320) );
  XOR U10138 ( .A(n10151), .B(n10323), .Z(n10144) );
  IV U10139 ( .A(n10150), .Z(n10323) );
  XNOR U10140 ( .A(n10147), .B(n10324), .Z(n10150) );
  XOR U10141 ( .A(n10325), .B(n10326), .Z(n10147) );
  ANDN U10142 ( .A(n10327), .B(n10328), .Z(n10326) );
  XNOR U10143 ( .A(n10325), .B(n10329), .Z(n10327) );
  XOR U10144 ( .A(n10158), .B(n10330), .Z(n10151) );
  IV U10145 ( .A(n10157), .Z(n10330) );
  XNOR U10146 ( .A(n10154), .B(n10331), .Z(n10157) );
  XOR U10147 ( .A(n10332), .B(n10333), .Z(n10154) );
  ANDN U10148 ( .A(n10334), .B(n10335), .Z(n10333) );
  XNOR U10149 ( .A(n10332), .B(n10336), .Z(n10334) );
  XOR U10150 ( .A(n10165), .B(n10337), .Z(n10158) );
  IV U10151 ( .A(n10164), .Z(n10337) );
  XNOR U10152 ( .A(n10161), .B(n10338), .Z(n10164) );
  XOR U10153 ( .A(n10339), .B(n10340), .Z(n10161) );
  ANDN U10154 ( .A(n10341), .B(n10342), .Z(n10340) );
  XNOR U10155 ( .A(n10339), .B(n10343), .Z(n10341) );
  XOR U10156 ( .A(n10172), .B(n10344), .Z(n10165) );
  IV U10157 ( .A(n10171), .Z(n10344) );
  XNOR U10158 ( .A(n10168), .B(n10345), .Z(n10171) );
  XOR U10159 ( .A(n10346), .B(n10347), .Z(n10168) );
  ANDN U10160 ( .A(n10348), .B(n10349), .Z(n10347) );
  XNOR U10161 ( .A(n10346), .B(n10350), .Z(n10348) );
  XOR U10162 ( .A(n10179), .B(n10351), .Z(n10172) );
  IV U10163 ( .A(n10178), .Z(n10351) );
  XNOR U10164 ( .A(n10175), .B(n10352), .Z(n10178) );
  XOR U10165 ( .A(n10353), .B(n10354), .Z(n10175) );
  ANDN U10166 ( .A(n10355), .B(n10356), .Z(n10354) );
  XNOR U10167 ( .A(n10353), .B(n10357), .Z(n10355) );
  XOR U10168 ( .A(n10186), .B(n10358), .Z(n10179) );
  IV U10169 ( .A(n10185), .Z(n10358) );
  XNOR U10170 ( .A(n10182), .B(n10359), .Z(n10185) );
  XOR U10171 ( .A(n10360), .B(n10361), .Z(n10182) );
  ANDN U10172 ( .A(n10362), .B(n10363), .Z(n10361) );
  XNOR U10173 ( .A(n10360), .B(n10364), .Z(n10362) );
  XOR U10174 ( .A(n10193), .B(n10365), .Z(n10186) );
  IV U10175 ( .A(n10192), .Z(n10365) );
  XNOR U10176 ( .A(n10189), .B(n10366), .Z(n10192) );
  XOR U10177 ( .A(n10367), .B(n10368), .Z(n10189) );
  ANDN U10178 ( .A(n10369), .B(n10370), .Z(n10368) );
  XNOR U10179 ( .A(n10367), .B(n10371), .Z(n10369) );
  XOR U10180 ( .A(n10200), .B(n10372), .Z(n10193) );
  IV U10181 ( .A(n10199), .Z(n10372) );
  XNOR U10182 ( .A(n10196), .B(n10373), .Z(n10199) );
  XOR U10183 ( .A(n10374), .B(n10375), .Z(n10196) );
  ANDN U10184 ( .A(n10376), .B(n10377), .Z(n10375) );
  XNOR U10185 ( .A(n10374), .B(n10378), .Z(n10376) );
  XOR U10186 ( .A(n10207), .B(n10379), .Z(n10200) );
  IV U10187 ( .A(n10206), .Z(n10379) );
  XNOR U10188 ( .A(n10203), .B(n10380), .Z(n10206) );
  XOR U10189 ( .A(n10381), .B(n10382), .Z(n10203) );
  ANDN U10190 ( .A(n10383), .B(n10384), .Z(n10382) );
  XNOR U10191 ( .A(n10381), .B(n10385), .Z(n10383) );
  XOR U10192 ( .A(n10213), .B(n10386), .Z(n10207) );
  IV U10193 ( .A(n10212), .Z(n10386) );
  XNOR U10194 ( .A(n10209), .B(n10387), .Z(n10212) );
  XOR U10195 ( .A(n10388), .B(n10389), .Z(n10209) );
  ANDN U10196 ( .A(n10390), .B(n10391), .Z(n10389) );
  XNOR U10197 ( .A(n10388), .B(n10392), .Z(n10390) );
  XOR U10198 ( .A(n10219), .B(n10393), .Z(n10213) );
  IV U10199 ( .A(n10218), .Z(n10393) );
  XNOR U10200 ( .A(n10215), .B(n10380), .Z(n10218) );
  AND U10201 ( .A(n10731), .B(n10017), .Z(n10380) );
  XOR U10202 ( .A(n10394), .B(n10395), .Z(n10215) );
  ANDN U10203 ( .A(n10396), .B(n10397), .Z(n10395) );
  XNOR U10204 ( .A(n10394), .B(n10398), .Z(n10396) );
  XOR U10205 ( .A(n10225), .B(n10399), .Z(n10219) );
  IV U10206 ( .A(n10224), .Z(n10399) );
  XNOR U10207 ( .A(n10221), .B(n10373), .Z(n10224) );
  AND U10208 ( .A(n11049), .B(n9621), .Z(n10373) );
  XOR U10209 ( .A(n10400), .B(n10401), .Z(n10221) );
  ANDN U10210 ( .A(n10402), .B(n10403), .Z(n10401) );
  XNOR U10211 ( .A(n10400), .B(n10404), .Z(n10402) );
  XOR U10212 ( .A(n10231), .B(n10405), .Z(n10225) );
  IV U10213 ( .A(n10230), .Z(n10405) );
  XNOR U10214 ( .A(n10227), .B(n10366), .Z(n10230) );
  AND U10215 ( .A(n11341), .B(n9198), .Z(n10366) );
  XOR U10216 ( .A(n10406), .B(n10407), .Z(n10227) );
  ANDN U10217 ( .A(n10408), .B(n10409), .Z(n10407) );
  XNOR U10218 ( .A(n10406), .B(n10410), .Z(n10408) );
  XOR U10219 ( .A(n10237), .B(n10411), .Z(n10231) );
  IV U10220 ( .A(n10236), .Z(n10411) );
  XNOR U10221 ( .A(n10233), .B(n10359), .Z(n10236) );
  AND U10222 ( .A(n11607), .B(n8748), .Z(n10359) );
  XOR U10223 ( .A(n10412), .B(n10413), .Z(n10233) );
  ANDN U10224 ( .A(n10414), .B(n10415), .Z(n10413) );
  XNOR U10225 ( .A(n10412), .B(n10416), .Z(n10414) );
  XOR U10226 ( .A(n10243), .B(n10417), .Z(n10237) );
  IV U10227 ( .A(n10242), .Z(n10417) );
  XNOR U10228 ( .A(n10239), .B(n10352), .Z(n10242) );
  AND U10229 ( .A(n11869), .B(n8272), .Z(n10352) );
  XOR U10230 ( .A(n10418), .B(n10419), .Z(n10239) );
  ANDN U10231 ( .A(n10420), .B(n10421), .Z(n10419) );
  XNOR U10232 ( .A(n10418), .B(n10422), .Z(n10420) );
  XOR U10233 ( .A(n10249), .B(n10423), .Z(n10243) );
  IV U10234 ( .A(n10248), .Z(n10423) );
  XNOR U10235 ( .A(n10245), .B(n10345), .Z(n10248) );
  AND U10236 ( .A(n12128), .B(n7770), .Z(n10345) );
  XOR U10237 ( .A(n10424), .B(n10425), .Z(n10245) );
  ANDN U10238 ( .A(n10426), .B(n10427), .Z(n10425) );
  XNOR U10239 ( .A(n10424), .B(n10428), .Z(n10426) );
  XOR U10240 ( .A(n10255), .B(n10429), .Z(n10249) );
  IV U10241 ( .A(n10254), .Z(n10429) );
  XNOR U10242 ( .A(n10251), .B(n10338), .Z(n10254) );
  AND U10243 ( .A(n12387), .B(n7241), .Z(n10338) );
  XOR U10244 ( .A(n10430), .B(n10431), .Z(n10251) );
  ANDN U10245 ( .A(n10432), .B(n10433), .Z(n10431) );
  XNOR U10246 ( .A(n10430), .B(n10434), .Z(n10432) );
  XOR U10247 ( .A(n10261), .B(n10435), .Z(n10255) );
  IV U10248 ( .A(n10260), .Z(n10435) );
  XNOR U10249 ( .A(n10257), .B(n10331), .Z(n10260) );
  AND U10250 ( .A(n12644), .B(n6688), .Z(n10331) );
  XOR U10251 ( .A(n10436), .B(n10437), .Z(n10257) );
  ANDN U10252 ( .A(n10438), .B(n10439), .Z(n10437) );
  XNOR U10253 ( .A(n10436), .B(n10440), .Z(n10438) );
  XOR U10254 ( .A(n10267), .B(n10441), .Z(n10261) );
  IV U10255 ( .A(n10266), .Z(n10441) );
  XNOR U10256 ( .A(n10263), .B(n10324), .Z(n10266) );
  AND U10257 ( .A(n12880), .B(n6118), .Z(n10324) );
  XOR U10258 ( .A(n10442), .B(n10443), .Z(n10263) );
  ANDN U10259 ( .A(n10444), .B(n10445), .Z(n10443) );
  XNOR U10260 ( .A(n10442), .B(n10446), .Z(n10444) );
  XOR U10261 ( .A(n10273), .B(n10447), .Z(n10267) );
  IV U10262 ( .A(n10272), .Z(n10447) );
  XNOR U10263 ( .A(n10269), .B(n10317), .Z(n10272) );
  AND U10264 ( .A(n13070), .B(n5561), .Z(n10317) );
  XOR U10265 ( .A(n10448), .B(n10449), .Z(n10269) );
  ANDN U10266 ( .A(n10450), .B(n10451), .Z(n10449) );
  XNOR U10267 ( .A(n10448), .B(n10452), .Z(n10450) );
  XOR U10268 ( .A(n10279), .B(n10453), .Z(n10273) );
  IV U10269 ( .A(n10278), .Z(n10453) );
  XNOR U10270 ( .A(n10275), .B(n10310), .Z(n10278) );
  AND U10271 ( .A(n13207), .B(n5030), .Z(n10310) );
  XOR U10272 ( .A(n10454), .B(n10455), .Z(n10275) );
  ANDN U10273 ( .A(n10456), .B(n10457), .Z(n10455) );
  XNOR U10274 ( .A(n10454), .B(n10458), .Z(n10456) );
  XNOR U10275 ( .A(n10284), .B(n10122), .Z(n10279) );
  XNOR U10276 ( .A(n10281), .B(n10459), .Z(n10284) );
  AND U10277 ( .A(n6527), .B(n4525), .Z(n10459) );
  XOR U10278 ( .A(n10460), .B(n10461), .Z(n10281) );
  ANDN U10279 ( .A(n10462), .B(n10463), .Z(n10461) );
  XNOR U10280 ( .A(n10307), .B(n10460), .Z(n10462) );
  XOR U10281 ( .A(n10464), .B(n10122), .Z(n10304) );
  NANDN U10282 ( .B(n6808), .A(n4046), .Z(n10122) );
  XOR U10283 ( .A(n10465), .B(n10466), .Z(n4046) );
  AND U10284 ( .A(n6809), .B(n10467), .Z(n10466) );
  XNOR U10285 ( .A(n10465), .B(n10291), .Z(n10467) );
  XOR U10286 ( .A(n10289), .B(n10465), .Z(n10291) );
  XOR U10287 ( .A(n10468), .B(n10469), .Z(n10289) );
  ANDN U10288 ( .A(n10468), .B(n10470), .Z(n10469) );
  XOR U10289 ( .A(n10471), .B(n7368), .Z(n10465) );
  IV U10290 ( .A(n10293), .Z(n10464) );
  XOR U10291 ( .A(n10472), .B(n10473), .Z(n10293) );
  AND U10292 ( .A(n10474), .B(n10475), .Z(n10473) );
  XNOR U10293 ( .A(n10476), .B(n10472), .Z(n10475) );
  XNOR U10294 ( .A(n10297), .B(n10300), .Z(n10303) );
  XOR U10295 ( .A(n10477), .B(n10478), .Z(n10297) );
  XOR U10296 ( .A(n10479), .B(n10480), .Z(n10300) );
  AND U10297 ( .A(n10479), .B(n10481), .Z(n10480) );
  XOR U10298 ( .A(n10482), .B(n10474), .Z(n10481) );
  XOR U10299 ( .A(n10483), .B(n10308), .Z(n10474) );
  XOR U10300 ( .A(n10315), .B(n10484), .Z(n10308) );
  IV U10301 ( .A(n10313), .Z(n10484) );
  XNOR U10302 ( .A(n10485), .B(n10312), .Z(n10313) );
  OR U10303 ( .A(n10486), .B(n10487), .Z(n10312) );
  NANDN U10304 ( .B(n6541), .A(n5030), .Z(n10485) );
  XOR U10305 ( .A(n10322), .B(n10488), .Z(n10315) );
  IV U10306 ( .A(n10321), .Z(n10488) );
  XNOR U10307 ( .A(n10318), .B(n10489), .Z(n10321) );
  XOR U10308 ( .A(n10490), .B(n10491), .Z(n10318) );
  NANDN U10309 ( .B(n10492), .A(n10493), .Z(n10490) );
  XOR U10310 ( .A(n10491), .B(n10494), .Z(n10493) );
  XOR U10311 ( .A(n10329), .B(n10495), .Z(n10322) );
  IV U10312 ( .A(n10328), .Z(n10495) );
  XNOR U10313 ( .A(n10325), .B(n10496), .Z(n10328) );
  XOR U10314 ( .A(n10497), .B(n10498), .Z(n10325) );
  ANDN U10315 ( .A(n10499), .B(n10500), .Z(n10498) );
  XNOR U10316 ( .A(n10497), .B(n10501), .Z(n10499) );
  XOR U10317 ( .A(n10336), .B(n10502), .Z(n10329) );
  IV U10318 ( .A(n10335), .Z(n10502) );
  XNOR U10319 ( .A(n10332), .B(n10503), .Z(n10335) );
  XOR U10320 ( .A(n10504), .B(n10505), .Z(n10332) );
  ANDN U10321 ( .A(n10506), .B(n10507), .Z(n10505) );
  XNOR U10322 ( .A(n10504), .B(n10508), .Z(n10506) );
  XOR U10323 ( .A(n10343), .B(n10509), .Z(n10336) );
  IV U10324 ( .A(n10342), .Z(n10509) );
  XNOR U10325 ( .A(n10339), .B(n10510), .Z(n10342) );
  XOR U10326 ( .A(n10511), .B(n10512), .Z(n10339) );
  ANDN U10327 ( .A(n10513), .B(n10514), .Z(n10512) );
  XNOR U10328 ( .A(n10511), .B(n10515), .Z(n10513) );
  XOR U10329 ( .A(n10350), .B(n10516), .Z(n10343) );
  IV U10330 ( .A(n10349), .Z(n10516) );
  XNOR U10331 ( .A(n10346), .B(n10517), .Z(n10349) );
  XOR U10332 ( .A(n10518), .B(n10519), .Z(n10346) );
  ANDN U10333 ( .A(n10520), .B(n10521), .Z(n10519) );
  XNOR U10334 ( .A(n10518), .B(n10522), .Z(n10520) );
  XOR U10335 ( .A(n10357), .B(n10523), .Z(n10350) );
  IV U10336 ( .A(n10356), .Z(n10523) );
  XNOR U10337 ( .A(n10353), .B(n10524), .Z(n10356) );
  XOR U10338 ( .A(n10525), .B(n10526), .Z(n10353) );
  ANDN U10339 ( .A(n10527), .B(n10528), .Z(n10526) );
  XNOR U10340 ( .A(n10525), .B(n10529), .Z(n10527) );
  XOR U10341 ( .A(n10364), .B(n10530), .Z(n10357) );
  IV U10342 ( .A(n10363), .Z(n10530) );
  XNOR U10343 ( .A(n10360), .B(n10531), .Z(n10363) );
  XOR U10344 ( .A(n10532), .B(n10533), .Z(n10360) );
  ANDN U10345 ( .A(n10534), .B(n10535), .Z(n10533) );
  XNOR U10346 ( .A(n10532), .B(n10536), .Z(n10534) );
  XOR U10347 ( .A(n10371), .B(n10537), .Z(n10364) );
  IV U10348 ( .A(n10370), .Z(n10537) );
  XNOR U10349 ( .A(n10367), .B(n10538), .Z(n10370) );
  XOR U10350 ( .A(n10539), .B(n10540), .Z(n10367) );
  ANDN U10351 ( .A(n10541), .B(n10542), .Z(n10540) );
  XNOR U10352 ( .A(n10539), .B(n10543), .Z(n10541) );
  XOR U10353 ( .A(n10378), .B(n10544), .Z(n10371) );
  IV U10354 ( .A(n10377), .Z(n10544) );
  XNOR U10355 ( .A(n10374), .B(n10545), .Z(n10377) );
  XOR U10356 ( .A(n10546), .B(n10547), .Z(n10374) );
  ANDN U10357 ( .A(n10548), .B(n10549), .Z(n10547) );
  XNOR U10358 ( .A(n10546), .B(n10550), .Z(n10548) );
  XOR U10359 ( .A(n10385), .B(n10551), .Z(n10378) );
  IV U10360 ( .A(n10384), .Z(n10551) );
  XNOR U10361 ( .A(n10381), .B(n10552), .Z(n10384) );
  XOR U10362 ( .A(n10553), .B(n10554), .Z(n10381) );
  ANDN U10363 ( .A(n10555), .B(n10556), .Z(n10554) );
  XNOR U10364 ( .A(n10553), .B(n10557), .Z(n10555) );
  XOR U10365 ( .A(n10392), .B(n10558), .Z(n10385) );
  IV U10366 ( .A(n10391), .Z(n10558) );
  XNOR U10367 ( .A(n10388), .B(n10559), .Z(n10391) );
  XOR U10368 ( .A(n10560), .B(n10561), .Z(n10388) );
  ANDN U10369 ( .A(n10562), .B(n10563), .Z(n10561) );
  XNOR U10370 ( .A(n10560), .B(n10564), .Z(n10562) );
  XOR U10371 ( .A(n10398), .B(n10565), .Z(n10392) );
  IV U10372 ( .A(n10397), .Z(n10565) );
  XNOR U10373 ( .A(n10394), .B(n10559), .Z(n10397) );
  AND U10374 ( .A(n10731), .B(n10387), .Z(n10559) );
  XOR U10375 ( .A(n10566), .B(n10567), .Z(n10394) );
  ANDN U10376 ( .A(n10568), .B(n10569), .Z(n10567) );
  XNOR U10377 ( .A(n10566), .B(n10570), .Z(n10568) );
  XOR U10378 ( .A(n10404), .B(n10571), .Z(n10398) );
  IV U10379 ( .A(n10403), .Z(n10571) );
  XNOR U10380 ( .A(n10400), .B(n10552), .Z(n10403) );
  AND U10381 ( .A(n11049), .B(n10017), .Z(n10552) );
  XOR U10382 ( .A(n10572), .B(n10573), .Z(n10400) );
  ANDN U10383 ( .A(n10574), .B(n10575), .Z(n10573) );
  XNOR U10384 ( .A(n10572), .B(n10576), .Z(n10574) );
  XOR U10385 ( .A(n10410), .B(n10577), .Z(n10404) );
  IV U10386 ( .A(n10409), .Z(n10577) );
  XNOR U10387 ( .A(n10406), .B(n10545), .Z(n10409) );
  AND U10388 ( .A(n11341), .B(n9621), .Z(n10545) );
  XOR U10389 ( .A(n10578), .B(n10579), .Z(n10406) );
  ANDN U10390 ( .A(n10580), .B(n10581), .Z(n10579) );
  XNOR U10391 ( .A(n10578), .B(n10582), .Z(n10580) );
  XOR U10392 ( .A(n10416), .B(n10583), .Z(n10410) );
  IV U10393 ( .A(n10415), .Z(n10583) );
  XNOR U10394 ( .A(n10412), .B(n10538), .Z(n10415) );
  AND U10395 ( .A(n11607), .B(n9198), .Z(n10538) );
  XOR U10396 ( .A(n10584), .B(n10585), .Z(n10412) );
  ANDN U10397 ( .A(n10586), .B(n10587), .Z(n10585) );
  XNOR U10398 ( .A(n10584), .B(n10588), .Z(n10586) );
  XOR U10399 ( .A(n10422), .B(n10589), .Z(n10416) );
  IV U10400 ( .A(n10421), .Z(n10589) );
  XNOR U10401 ( .A(n10418), .B(n10531), .Z(n10421) );
  AND U10402 ( .A(n11869), .B(n8748), .Z(n10531) );
  XOR U10403 ( .A(n10590), .B(n10591), .Z(n10418) );
  ANDN U10404 ( .A(n10592), .B(n10593), .Z(n10591) );
  XNOR U10405 ( .A(n10590), .B(n10594), .Z(n10592) );
  XOR U10406 ( .A(n10428), .B(n10595), .Z(n10422) );
  IV U10407 ( .A(n10427), .Z(n10595) );
  XNOR U10408 ( .A(n10424), .B(n10524), .Z(n10427) );
  AND U10409 ( .A(n12128), .B(n8272), .Z(n10524) );
  XOR U10410 ( .A(n10596), .B(n10597), .Z(n10424) );
  ANDN U10411 ( .A(n10598), .B(n10599), .Z(n10597) );
  XNOR U10412 ( .A(n10596), .B(n10600), .Z(n10598) );
  XOR U10413 ( .A(n10434), .B(n10601), .Z(n10428) );
  IV U10414 ( .A(n10433), .Z(n10601) );
  XNOR U10415 ( .A(n10430), .B(n10517), .Z(n10433) );
  AND U10416 ( .A(n12387), .B(n7770), .Z(n10517) );
  XOR U10417 ( .A(n10602), .B(n10603), .Z(n10430) );
  ANDN U10418 ( .A(n10604), .B(n10605), .Z(n10603) );
  XNOR U10419 ( .A(n10602), .B(n10606), .Z(n10604) );
  XOR U10420 ( .A(n10440), .B(n10607), .Z(n10434) );
  IV U10421 ( .A(n10439), .Z(n10607) );
  XNOR U10422 ( .A(n10436), .B(n10510), .Z(n10439) );
  AND U10423 ( .A(n12644), .B(n7241), .Z(n10510) );
  XOR U10424 ( .A(n10608), .B(n10609), .Z(n10436) );
  ANDN U10425 ( .A(n10610), .B(n10611), .Z(n10609) );
  XNOR U10426 ( .A(n10608), .B(n10612), .Z(n10610) );
  XOR U10427 ( .A(n10446), .B(n10613), .Z(n10440) );
  IV U10428 ( .A(n10445), .Z(n10613) );
  XNOR U10429 ( .A(n10442), .B(n10503), .Z(n10445) );
  AND U10430 ( .A(n12880), .B(n6688), .Z(n10503) );
  XOR U10431 ( .A(n10614), .B(n10615), .Z(n10442) );
  ANDN U10432 ( .A(n10616), .B(n10617), .Z(n10615) );
  XNOR U10433 ( .A(n10614), .B(n10618), .Z(n10616) );
  XOR U10434 ( .A(n10452), .B(n10619), .Z(n10446) );
  IV U10435 ( .A(n10451), .Z(n10619) );
  XNOR U10436 ( .A(n10448), .B(n10496), .Z(n10451) );
  AND U10437 ( .A(n13070), .B(n6118), .Z(n10496) );
  XOR U10438 ( .A(n10620), .B(n10621), .Z(n10448) );
  ANDN U10439 ( .A(n10622), .B(n10623), .Z(n10621) );
  XNOR U10440 ( .A(n10620), .B(n10624), .Z(n10622) );
  XOR U10441 ( .A(n10458), .B(n10625), .Z(n10452) );
  IV U10442 ( .A(n10457), .Z(n10625) );
  XNOR U10443 ( .A(n10454), .B(n10489), .Z(n10457) );
  AND U10444 ( .A(n13207), .B(n5561), .Z(n10489) );
  XOR U10445 ( .A(n10626), .B(n10627), .Z(n10454) );
  ANDN U10446 ( .A(n10628), .B(n10629), .Z(n10627) );
  XNOR U10447 ( .A(n10626), .B(n10630), .Z(n10628) );
  XNOR U10448 ( .A(n10463), .B(n10307), .Z(n10458) );
  XNOR U10449 ( .A(n10460), .B(n10631), .Z(n10463) );
  AND U10450 ( .A(n6527), .B(n5030), .Z(n10631) );
  XOR U10451 ( .A(n10632), .B(n10633), .Z(n10460) );
  ANDN U10452 ( .A(n10634), .B(n10635), .Z(n10633) );
  XNOR U10453 ( .A(n10486), .B(n10632), .Z(n10634) );
  XOR U10454 ( .A(n10636), .B(n10307), .Z(n10483) );
  NANDN U10455 ( .B(n6808), .A(n4525), .Z(n10307) );
  XOR U10456 ( .A(n10637), .B(n10638), .Z(n4525) );
  AND U10457 ( .A(n6809), .B(n10639), .Z(n10638) );
  XNOR U10458 ( .A(n10637), .B(n10470), .Z(n10639) );
  XOR U10459 ( .A(n10468), .B(n10637), .Z(n10470) );
  XOR U10460 ( .A(n10640), .B(n10641), .Z(n10468) );
  ANDN U10461 ( .A(n10640), .B(n10642), .Z(n10641) );
  XOR U10462 ( .A(n10643), .B(n7368), .Z(n10637) );
  IV U10463 ( .A(n10472), .Z(n10636) );
  XOR U10464 ( .A(n10644), .B(n10645), .Z(n10472) );
  AND U10465 ( .A(n10646), .B(n10647), .Z(n10645) );
  XNOR U10466 ( .A(n10648), .B(n10644), .Z(n10647) );
  XNOR U10467 ( .A(n10476), .B(n10479), .Z(n10482) );
  XOR U10468 ( .A(n10649), .B(n10650), .Z(n10476) );
  XOR U10469 ( .A(n10651), .B(n10652), .Z(n10479) );
  AND U10470 ( .A(n10651), .B(n10653), .Z(n10652) );
  XOR U10471 ( .A(n10654), .B(n10646), .Z(n10653) );
  XOR U10472 ( .A(n10655), .B(n10487), .Z(n10646) );
  XOR U10473 ( .A(n10494), .B(n10656), .Z(n10487) );
  IV U10474 ( .A(n10492), .Z(n10656) );
  XNOR U10475 ( .A(n10657), .B(n10491), .Z(n10492) );
  OR U10476 ( .A(n10658), .B(n10659), .Z(n10491) );
  NANDN U10477 ( .B(n6541), .A(n5561), .Z(n10657) );
  XOR U10478 ( .A(n10501), .B(n10660), .Z(n10494) );
  IV U10479 ( .A(n10500), .Z(n10660) );
  XNOR U10480 ( .A(n10497), .B(n10661), .Z(n10500) );
  XOR U10481 ( .A(n10662), .B(n10663), .Z(n10497) );
  NANDN U10482 ( .B(n10664), .A(n10665), .Z(n10662) );
  XOR U10483 ( .A(n10663), .B(n10666), .Z(n10665) );
  XOR U10484 ( .A(n10508), .B(n10667), .Z(n10501) );
  IV U10485 ( .A(n10507), .Z(n10667) );
  XNOR U10486 ( .A(n10504), .B(n10668), .Z(n10507) );
  XOR U10487 ( .A(n10669), .B(n10670), .Z(n10504) );
  ANDN U10488 ( .A(n10671), .B(n10672), .Z(n10670) );
  XNOR U10489 ( .A(n10669), .B(n10673), .Z(n10671) );
  XOR U10490 ( .A(n10515), .B(n10674), .Z(n10508) );
  IV U10491 ( .A(n10514), .Z(n10674) );
  XNOR U10492 ( .A(n10511), .B(n10675), .Z(n10514) );
  XOR U10493 ( .A(n10676), .B(n10677), .Z(n10511) );
  ANDN U10494 ( .A(n10678), .B(n10679), .Z(n10677) );
  XNOR U10495 ( .A(n10676), .B(n10680), .Z(n10678) );
  XOR U10496 ( .A(n10522), .B(n10681), .Z(n10515) );
  IV U10497 ( .A(n10521), .Z(n10681) );
  XNOR U10498 ( .A(n10518), .B(n10682), .Z(n10521) );
  XOR U10499 ( .A(n10683), .B(n10684), .Z(n10518) );
  ANDN U10500 ( .A(n10685), .B(n10686), .Z(n10684) );
  XNOR U10501 ( .A(n10683), .B(n10687), .Z(n10685) );
  XOR U10502 ( .A(n10529), .B(n10688), .Z(n10522) );
  IV U10503 ( .A(n10528), .Z(n10688) );
  XNOR U10504 ( .A(n10525), .B(n10689), .Z(n10528) );
  XOR U10505 ( .A(n10690), .B(n10691), .Z(n10525) );
  ANDN U10506 ( .A(n10692), .B(n10693), .Z(n10691) );
  XNOR U10507 ( .A(n10690), .B(n10694), .Z(n10692) );
  XOR U10508 ( .A(n10536), .B(n10695), .Z(n10529) );
  IV U10509 ( .A(n10535), .Z(n10695) );
  XNOR U10510 ( .A(n10532), .B(n10696), .Z(n10535) );
  XOR U10511 ( .A(n10697), .B(n10698), .Z(n10532) );
  ANDN U10512 ( .A(n10699), .B(n10700), .Z(n10698) );
  XNOR U10513 ( .A(n10697), .B(n10701), .Z(n10699) );
  XOR U10514 ( .A(n10543), .B(n10702), .Z(n10536) );
  IV U10515 ( .A(n10542), .Z(n10702) );
  XNOR U10516 ( .A(n10539), .B(n10703), .Z(n10542) );
  XOR U10517 ( .A(n10704), .B(n10705), .Z(n10539) );
  ANDN U10518 ( .A(n10706), .B(n10707), .Z(n10705) );
  XNOR U10519 ( .A(n10704), .B(n10708), .Z(n10706) );
  XOR U10520 ( .A(n10550), .B(n10709), .Z(n10543) );
  IV U10521 ( .A(n10549), .Z(n10709) );
  XNOR U10522 ( .A(n10546), .B(n10710), .Z(n10549) );
  XOR U10523 ( .A(n10711), .B(n10712), .Z(n10546) );
  ANDN U10524 ( .A(n10713), .B(n10714), .Z(n10712) );
  XNOR U10525 ( .A(n10711), .B(n10715), .Z(n10713) );
  XOR U10526 ( .A(n10557), .B(n10716), .Z(n10550) );
  IV U10527 ( .A(n10556), .Z(n10716) );
  XNOR U10528 ( .A(n10553), .B(n10717), .Z(n10556) );
  XOR U10529 ( .A(n10718), .B(n10719), .Z(n10553) );
  ANDN U10530 ( .A(n10720), .B(n10721), .Z(n10719) );
  XNOR U10531 ( .A(n10718), .B(n10722), .Z(n10720) );
  XOR U10532 ( .A(n10564), .B(n10723), .Z(n10557) );
  IV U10533 ( .A(n10563), .Z(n10723) );
  XNOR U10534 ( .A(n10560), .B(n10724), .Z(n10563) );
  XOR U10535 ( .A(n10725), .B(n10726), .Z(n10560) );
  ANDN U10536 ( .A(n10727), .B(n10728), .Z(n10726) );
  XNOR U10537 ( .A(n10725), .B(n10729), .Z(n10727) );
  XOR U10538 ( .A(n10570), .B(n10730), .Z(n10564) );
  IV U10539 ( .A(n10569), .Z(n10730) );
  XNOR U10540 ( .A(n10566), .B(n10731), .Z(n10569) );
  XOR U10541 ( .A(n10732), .B(n10733), .Z(n10566) );
  ANDN U10542 ( .A(n10734), .B(n10735), .Z(n10733) );
  XNOR U10543 ( .A(n10732), .B(n10736), .Z(n10734) );
  XOR U10544 ( .A(n10576), .B(n10737), .Z(n10570) );
  IV U10545 ( .A(n10575), .Z(n10737) );
  XNOR U10546 ( .A(n10572), .B(n10724), .Z(n10575) );
  AND U10547 ( .A(n11049), .B(n10387), .Z(n10724) );
  XOR U10548 ( .A(n10738), .B(n10739), .Z(n10572) );
  ANDN U10549 ( .A(n10740), .B(n10741), .Z(n10739) );
  XNOR U10550 ( .A(n10738), .B(n10742), .Z(n10740) );
  XOR U10551 ( .A(n10582), .B(n10743), .Z(n10576) );
  IV U10552 ( .A(n10581), .Z(n10743) );
  XNOR U10553 ( .A(n10578), .B(n10717), .Z(n10581) );
  AND U10554 ( .A(n11341), .B(n10017), .Z(n10717) );
  XOR U10555 ( .A(n10744), .B(n10745), .Z(n10578) );
  ANDN U10556 ( .A(n10746), .B(n10747), .Z(n10745) );
  XNOR U10557 ( .A(n10744), .B(n10748), .Z(n10746) );
  XOR U10558 ( .A(n10588), .B(n10749), .Z(n10582) );
  IV U10559 ( .A(n10587), .Z(n10749) );
  XNOR U10560 ( .A(n10584), .B(n10710), .Z(n10587) );
  AND U10561 ( .A(n11607), .B(n9621), .Z(n10710) );
  XOR U10562 ( .A(n10750), .B(n10751), .Z(n10584) );
  ANDN U10563 ( .A(n10752), .B(n10753), .Z(n10751) );
  XNOR U10564 ( .A(n10750), .B(n10754), .Z(n10752) );
  XOR U10565 ( .A(n10594), .B(n10755), .Z(n10588) );
  IV U10566 ( .A(n10593), .Z(n10755) );
  XNOR U10567 ( .A(n10590), .B(n10703), .Z(n10593) );
  AND U10568 ( .A(n11869), .B(n9198), .Z(n10703) );
  XOR U10569 ( .A(n10756), .B(n10757), .Z(n10590) );
  ANDN U10570 ( .A(n10758), .B(n10759), .Z(n10757) );
  XNOR U10571 ( .A(n10756), .B(n10760), .Z(n10758) );
  XOR U10572 ( .A(n10600), .B(n10761), .Z(n10594) );
  IV U10573 ( .A(n10599), .Z(n10761) );
  XNOR U10574 ( .A(n10596), .B(n10696), .Z(n10599) );
  AND U10575 ( .A(n12128), .B(n8748), .Z(n10696) );
  XOR U10576 ( .A(n10762), .B(n10763), .Z(n10596) );
  ANDN U10577 ( .A(n10764), .B(n10765), .Z(n10763) );
  XNOR U10578 ( .A(n10762), .B(n10766), .Z(n10764) );
  XOR U10579 ( .A(n10606), .B(n10767), .Z(n10600) );
  IV U10580 ( .A(n10605), .Z(n10767) );
  XNOR U10581 ( .A(n10602), .B(n10689), .Z(n10605) );
  AND U10582 ( .A(n12387), .B(n8272), .Z(n10689) );
  XOR U10583 ( .A(n10768), .B(n10769), .Z(n10602) );
  ANDN U10584 ( .A(n10770), .B(n10771), .Z(n10769) );
  XNOR U10585 ( .A(n10768), .B(n10772), .Z(n10770) );
  XOR U10586 ( .A(n10612), .B(n10773), .Z(n10606) );
  IV U10587 ( .A(n10611), .Z(n10773) );
  XNOR U10588 ( .A(n10608), .B(n10682), .Z(n10611) );
  AND U10589 ( .A(n12644), .B(n7770), .Z(n10682) );
  XOR U10590 ( .A(n10774), .B(n10775), .Z(n10608) );
  ANDN U10591 ( .A(n10776), .B(n10777), .Z(n10775) );
  XNOR U10592 ( .A(n10774), .B(n10778), .Z(n10776) );
  XOR U10593 ( .A(n10618), .B(n10779), .Z(n10612) );
  IV U10594 ( .A(n10617), .Z(n10779) );
  XNOR U10595 ( .A(n10614), .B(n10675), .Z(n10617) );
  AND U10596 ( .A(n12880), .B(n7241), .Z(n10675) );
  XOR U10597 ( .A(n10780), .B(n10781), .Z(n10614) );
  ANDN U10598 ( .A(n10782), .B(n10783), .Z(n10781) );
  XNOR U10599 ( .A(n10780), .B(n10784), .Z(n10782) );
  XOR U10600 ( .A(n10624), .B(n10785), .Z(n10618) );
  IV U10601 ( .A(n10623), .Z(n10785) );
  XNOR U10602 ( .A(n10620), .B(n10668), .Z(n10623) );
  AND U10603 ( .A(n13070), .B(n6688), .Z(n10668) );
  XOR U10604 ( .A(n10786), .B(n10787), .Z(n10620) );
  ANDN U10605 ( .A(n10788), .B(n10789), .Z(n10787) );
  XNOR U10606 ( .A(n10786), .B(n10790), .Z(n10788) );
  XOR U10607 ( .A(n10630), .B(n10791), .Z(n10624) );
  IV U10608 ( .A(n10629), .Z(n10791) );
  XNOR U10609 ( .A(n10626), .B(n10661), .Z(n10629) );
  AND U10610 ( .A(n13207), .B(n6118), .Z(n10661) );
  XOR U10611 ( .A(n10792), .B(n10793), .Z(n10626) );
  ANDN U10612 ( .A(n10794), .B(n10795), .Z(n10793) );
  XNOR U10613 ( .A(n10792), .B(n10796), .Z(n10794) );
  XNOR U10614 ( .A(n10635), .B(n10486), .Z(n10630) );
  XNOR U10615 ( .A(n10632), .B(n10797), .Z(n10635) );
  AND U10616 ( .A(n6527), .B(n5561), .Z(n10797) );
  XOR U10617 ( .A(n10798), .B(n10799), .Z(n10632) );
  ANDN U10618 ( .A(n10800), .B(n10801), .Z(n10799) );
  XNOR U10619 ( .A(n10658), .B(n10798), .Z(n10800) );
  XOR U10620 ( .A(n10802), .B(n10486), .Z(n10655) );
  NANDN U10621 ( .B(n6808), .A(n5030), .Z(n10486) );
  XOR U10622 ( .A(n10803), .B(n10804), .Z(n5030) );
  AND U10623 ( .A(n6809), .B(n10805), .Z(n10804) );
  XNOR U10624 ( .A(n10803), .B(n10642), .Z(n10805) );
  XOR U10625 ( .A(n10640), .B(n10803), .Z(n10642) );
  XOR U10626 ( .A(n10806), .B(n10807), .Z(n10640) );
  ANDN U10627 ( .A(n10806), .B(n10808), .Z(n10807) );
  XOR U10628 ( .A(n10809), .B(n7368), .Z(n10803) );
  IV U10629 ( .A(n10644), .Z(n10802) );
  XOR U10630 ( .A(n10810), .B(n10811), .Z(n10644) );
  AND U10631 ( .A(n10812), .B(n10813), .Z(n10811) );
  XNOR U10632 ( .A(n10814), .B(n10810), .Z(n10813) );
  XNOR U10633 ( .A(n10648), .B(n10651), .Z(n10654) );
  XOR U10634 ( .A(n10815), .B(n10816), .Z(n10648) );
  XOR U10635 ( .A(n10817), .B(n10818), .Z(n10651) );
  AND U10636 ( .A(n10817), .B(n10819), .Z(n10818) );
  XOR U10637 ( .A(n10820), .B(n10812), .Z(n10819) );
  XOR U10638 ( .A(n10821), .B(n10659), .Z(n10812) );
  XOR U10639 ( .A(n10666), .B(n10822), .Z(n10659) );
  IV U10640 ( .A(n10664), .Z(n10822) );
  XNOR U10641 ( .A(n10823), .B(n10663), .Z(n10664) );
  OR U10642 ( .A(n10824), .B(n10825), .Z(n10663) );
  NANDN U10643 ( .B(n6541), .A(n6118), .Z(n10823) );
  XOR U10644 ( .A(n10673), .B(n10826), .Z(n10666) );
  IV U10645 ( .A(n10672), .Z(n10826) );
  XNOR U10646 ( .A(n10669), .B(n10827), .Z(n10672) );
  XOR U10647 ( .A(n10828), .B(n10829), .Z(n10669) );
  NANDN U10648 ( .B(n10830), .A(n10831), .Z(n10828) );
  XOR U10649 ( .A(n10829), .B(n10832), .Z(n10831) );
  XOR U10650 ( .A(n10680), .B(n10833), .Z(n10673) );
  IV U10651 ( .A(n10679), .Z(n10833) );
  XNOR U10652 ( .A(n10676), .B(n10834), .Z(n10679) );
  XOR U10653 ( .A(n10835), .B(n10836), .Z(n10676) );
  ANDN U10654 ( .A(n10837), .B(n10838), .Z(n10836) );
  XNOR U10655 ( .A(n10835), .B(n10839), .Z(n10837) );
  XOR U10656 ( .A(n10687), .B(n10840), .Z(n10680) );
  IV U10657 ( .A(n10686), .Z(n10840) );
  XNOR U10658 ( .A(n10683), .B(n10841), .Z(n10686) );
  XOR U10659 ( .A(n10842), .B(n10843), .Z(n10683) );
  ANDN U10660 ( .A(n10844), .B(n10845), .Z(n10843) );
  XNOR U10661 ( .A(n10842), .B(n10846), .Z(n10844) );
  XOR U10662 ( .A(n10694), .B(n10847), .Z(n10687) );
  IV U10663 ( .A(n10693), .Z(n10847) );
  XNOR U10664 ( .A(n10690), .B(n10848), .Z(n10693) );
  XOR U10665 ( .A(n10849), .B(n10850), .Z(n10690) );
  ANDN U10666 ( .A(n10851), .B(n10852), .Z(n10850) );
  XNOR U10667 ( .A(n10849), .B(n10853), .Z(n10851) );
  XOR U10668 ( .A(n10701), .B(n10854), .Z(n10694) );
  IV U10669 ( .A(n10700), .Z(n10854) );
  XNOR U10670 ( .A(n10697), .B(n10855), .Z(n10700) );
  XOR U10671 ( .A(n10856), .B(n10857), .Z(n10697) );
  ANDN U10672 ( .A(n10858), .B(n10859), .Z(n10857) );
  XNOR U10673 ( .A(n10856), .B(n10860), .Z(n10858) );
  XOR U10674 ( .A(n10708), .B(n10861), .Z(n10701) );
  IV U10675 ( .A(n10707), .Z(n10861) );
  XNOR U10676 ( .A(n10704), .B(n10862), .Z(n10707) );
  XOR U10677 ( .A(n10863), .B(n10864), .Z(n10704) );
  ANDN U10678 ( .A(n10865), .B(n10866), .Z(n10864) );
  XNOR U10679 ( .A(n10863), .B(n10867), .Z(n10865) );
  XOR U10680 ( .A(n10715), .B(n10868), .Z(n10708) );
  IV U10681 ( .A(n10714), .Z(n10868) );
  XNOR U10682 ( .A(n10711), .B(n10869), .Z(n10714) );
  XOR U10683 ( .A(n10870), .B(n10871), .Z(n10711) );
  ANDN U10684 ( .A(n10872), .B(n10873), .Z(n10871) );
  XNOR U10685 ( .A(n10870), .B(n10874), .Z(n10872) );
  XOR U10686 ( .A(n10722), .B(n10875), .Z(n10715) );
  IV U10687 ( .A(n10721), .Z(n10875) );
  XNOR U10688 ( .A(n10718), .B(n10876), .Z(n10721) );
  XOR U10689 ( .A(n10877), .B(n10878), .Z(n10718) );
  ANDN U10690 ( .A(n10879), .B(n10880), .Z(n10878) );
  XNOR U10691 ( .A(n10877), .B(n10881), .Z(n10879) );
  XOR U10692 ( .A(n10729), .B(n10882), .Z(n10722) );
  IV U10693 ( .A(n10728), .Z(n10882) );
  XNOR U10694 ( .A(n10725), .B(n10883), .Z(n10728) );
  XOR U10695 ( .A(n10884), .B(n10885), .Z(n10725) );
  ANDN U10696 ( .A(n10886), .B(n10887), .Z(n10885) );
  XNOR U10697 ( .A(n10884), .B(n10888), .Z(n10886) );
  XOR U10698 ( .A(n10736), .B(n10889), .Z(n10729) );
  IV U10699 ( .A(n10735), .Z(n10889) );
  XNOR U10700 ( .A(n10732), .B(n10890), .Z(n10735) );
  XOR U10701 ( .A(n10891), .B(n10892), .Z(n10732) );
  ANDN U10702 ( .A(n10893), .B(n10894), .Z(n10892) );
  XNOR U10703 ( .A(n10891), .B(n10895), .Z(n10893) );
  XOR U10704 ( .A(n10742), .B(n10896), .Z(n10736) );
  IV U10705 ( .A(n10741), .Z(n10896) );
  XNOR U10706 ( .A(n10738), .B(n10890), .Z(n10741) );
  AND U10707 ( .A(n11049), .B(n10731), .Z(n10890) );
  XOR U10708 ( .A(n10897), .B(n10898), .Z(n10738) );
  ANDN U10709 ( .A(n10899), .B(n10900), .Z(n10898) );
  XNOR U10710 ( .A(n10897), .B(n10901), .Z(n10899) );
  XOR U10711 ( .A(n10748), .B(n10902), .Z(n10742) );
  IV U10712 ( .A(n10747), .Z(n10902) );
  XNOR U10713 ( .A(n10744), .B(n10883), .Z(n10747) );
  AND U10714 ( .A(n11341), .B(n10387), .Z(n10883) );
  XOR U10715 ( .A(n10903), .B(n10904), .Z(n10744) );
  ANDN U10716 ( .A(n10905), .B(n10906), .Z(n10904) );
  XNOR U10717 ( .A(n10903), .B(n10907), .Z(n10905) );
  XOR U10718 ( .A(n10754), .B(n10908), .Z(n10748) );
  IV U10719 ( .A(n10753), .Z(n10908) );
  XNOR U10720 ( .A(n10750), .B(n10876), .Z(n10753) );
  AND U10721 ( .A(n11607), .B(n10017), .Z(n10876) );
  XOR U10722 ( .A(n10909), .B(n10910), .Z(n10750) );
  ANDN U10723 ( .A(n10911), .B(n10912), .Z(n10910) );
  XNOR U10724 ( .A(n10909), .B(n10913), .Z(n10911) );
  XOR U10725 ( .A(n10760), .B(n10914), .Z(n10754) );
  IV U10726 ( .A(n10759), .Z(n10914) );
  XNOR U10727 ( .A(n10756), .B(n10869), .Z(n10759) );
  AND U10728 ( .A(n11869), .B(n9621), .Z(n10869) );
  XOR U10729 ( .A(n10915), .B(n10916), .Z(n10756) );
  ANDN U10730 ( .A(n10917), .B(n10918), .Z(n10916) );
  XNOR U10731 ( .A(n10915), .B(n10919), .Z(n10917) );
  XOR U10732 ( .A(n10766), .B(n10920), .Z(n10760) );
  IV U10733 ( .A(n10765), .Z(n10920) );
  XNOR U10734 ( .A(n10762), .B(n10862), .Z(n10765) );
  AND U10735 ( .A(n12128), .B(n9198), .Z(n10862) );
  XOR U10736 ( .A(n10921), .B(n10922), .Z(n10762) );
  ANDN U10737 ( .A(n10923), .B(n10924), .Z(n10922) );
  XNOR U10738 ( .A(n10921), .B(n10925), .Z(n10923) );
  XOR U10739 ( .A(n10772), .B(n10926), .Z(n10766) );
  IV U10740 ( .A(n10771), .Z(n10926) );
  XNOR U10741 ( .A(n10768), .B(n10855), .Z(n10771) );
  AND U10742 ( .A(n12387), .B(n8748), .Z(n10855) );
  XOR U10743 ( .A(n10927), .B(n10928), .Z(n10768) );
  ANDN U10744 ( .A(n10929), .B(n10930), .Z(n10928) );
  XNOR U10745 ( .A(n10927), .B(n10931), .Z(n10929) );
  XOR U10746 ( .A(n10778), .B(n10932), .Z(n10772) );
  IV U10747 ( .A(n10777), .Z(n10932) );
  XNOR U10748 ( .A(n10774), .B(n10848), .Z(n10777) );
  AND U10749 ( .A(n12644), .B(n8272), .Z(n10848) );
  XOR U10750 ( .A(n10933), .B(n10934), .Z(n10774) );
  ANDN U10751 ( .A(n10935), .B(n10936), .Z(n10934) );
  XNOR U10752 ( .A(n10933), .B(n10937), .Z(n10935) );
  XOR U10753 ( .A(n10784), .B(n10938), .Z(n10778) );
  IV U10754 ( .A(n10783), .Z(n10938) );
  XNOR U10755 ( .A(n10780), .B(n10841), .Z(n10783) );
  AND U10756 ( .A(n12880), .B(n7770), .Z(n10841) );
  XOR U10757 ( .A(n10939), .B(n10940), .Z(n10780) );
  ANDN U10758 ( .A(n10941), .B(n10942), .Z(n10940) );
  XNOR U10759 ( .A(n10939), .B(n10943), .Z(n10941) );
  XOR U10760 ( .A(n10790), .B(n10944), .Z(n10784) );
  IV U10761 ( .A(n10789), .Z(n10944) );
  XNOR U10762 ( .A(n10786), .B(n10834), .Z(n10789) );
  AND U10763 ( .A(n13070), .B(n7241), .Z(n10834) );
  XOR U10764 ( .A(n10945), .B(n10946), .Z(n10786) );
  ANDN U10765 ( .A(n10947), .B(n10948), .Z(n10946) );
  XNOR U10766 ( .A(n10945), .B(n10949), .Z(n10947) );
  XOR U10767 ( .A(n10796), .B(n10950), .Z(n10790) );
  IV U10768 ( .A(n10795), .Z(n10950) );
  XNOR U10769 ( .A(n10792), .B(n10827), .Z(n10795) );
  AND U10770 ( .A(n13207), .B(n6688), .Z(n10827) );
  XOR U10771 ( .A(n10951), .B(n10952), .Z(n10792) );
  ANDN U10772 ( .A(n10953), .B(n10954), .Z(n10952) );
  XNOR U10773 ( .A(n10951), .B(n10955), .Z(n10953) );
  XNOR U10774 ( .A(n10801), .B(n10658), .Z(n10796) );
  XNOR U10775 ( .A(n10798), .B(n10956), .Z(n10801) );
  AND U10776 ( .A(n6527), .B(n6118), .Z(n10956) );
  XOR U10777 ( .A(n10957), .B(n10958), .Z(n10798) );
  ANDN U10778 ( .A(n10959), .B(n10960), .Z(n10958) );
  XNOR U10779 ( .A(n10824), .B(n10957), .Z(n10959) );
  XOR U10780 ( .A(n10961), .B(n10658), .Z(n10821) );
  NANDN U10781 ( .B(n6808), .A(n5561), .Z(n10658) );
  XOR U10782 ( .A(n10962), .B(n10963), .Z(n5561) );
  AND U10783 ( .A(n6809), .B(n10964), .Z(n10963) );
  XNOR U10784 ( .A(n10962), .B(n10808), .Z(n10964) );
  XOR U10785 ( .A(n10806), .B(n10962), .Z(n10808) );
  XOR U10786 ( .A(n10965), .B(n10966), .Z(n10806) );
  ANDN U10787 ( .A(n10965), .B(n10967), .Z(n10966) );
  XOR U10788 ( .A(n10968), .B(n7368), .Z(n10962) );
  IV U10789 ( .A(n10810), .Z(n10961) );
  XOR U10790 ( .A(n10969), .B(n10970), .Z(n10810) );
  AND U10791 ( .A(n10971), .B(n10972), .Z(n10970) );
  XNOR U10792 ( .A(n10973), .B(n10969), .Z(n10972) );
  XNOR U10793 ( .A(n10814), .B(n10817), .Z(n10820) );
  XOR U10794 ( .A(n10974), .B(n10975), .Z(n10814) );
  XOR U10795 ( .A(n10976), .B(n10977), .Z(n10817) );
  AND U10796 ( .A(n10976), .B(n10978), .Z(n10977) );
  XOR U10797 ( .A(n10979), .B(n10971), .Z(n10978) );
  XOR U10798 ( .A(n10980), .B(n10825), .Z(n10971) );
  XOR U10799 ( .A(n10832), .B(n10981), .Z(n10825) );
  IV U10800 ( .A(n10830), .Z(n10981) );
  XNOR U10801 ( .A(n10982), .B(n10829), .Z(n10830) );
  OR U10802 ( .A(n10983), .B(n10984), .Z(n10829) );
  NANDN U10803 ( .B(n6541), .A(n6688), .Z(n10982) );
  XOR U10804 ( .A(n10839), .B(n10985), .Z(n10832) );
  IV U10805 ( .A(n10838), .Z(n10985) );
  XNOR U10806 ( .A(n10835), .B(n10986), .Z(n10838) );
  XOR U10807 ( .A(n10987), .B(n10988), .Z(n10835) );
  NANDN U10808 ( .B(n10989), .A(n10990), .Z(n10987) );
  XOR U10809 ( .A(n10988), .B(n10991), .Z(n10990) );
  XOR U10810 ( .A(n10846), .B(n10992), .Z(n10839) );
  IV U10811 ( .A(n10845), .Z(n10992) );
  XNOR U10812 ( .A(n10842), .B(n10993), .Z(n10845) );
  XOR U10813 ( .A(n10994), .B(n10995), .Z(n10842) );
  ANDN U10814 ( .A(n10996), .B(n10997), .Z(n10995) );
  XNOR U10815 ( .A(n10994), .B(n10998), .Z(n10996) );
  XOR U10816 ( .A(n10853), .B(n10999), .Z(n10846) );
  IV U10817 ( .A(n10852), .Z(n10999) );
  XNOR U10818 ( .A(n10849), .B(n11000), .Z(n10852) );
  XOR U10819 ( .A(n11001), .B(n11002), .Z(n10849) );
  ANDN U10820 ( .A(n11003), .B(n11004), .Z(n11002) );
  XNOR U10821 ( .A(n11001), .B(n11005), .Z(n11003) );
  XOR U10822 ( .A(n10860), .B(n11006), .Z(n10853) );
  IV U10823 ( .A(n10859), .Z(n11006) );
  XNOR U10824 ( .A(n10856), .B(n11007), .Z(n10859) );
  XOR U10825 ( .A(n11008), .B(n11009), .Z(n10856) );
  ANDN U10826 ( .A(n11010), .B(n11011), .Z(n11009) );
  XNOR U10827 ( .A(n11008), .B(n11012), .Z(n11010) );
  XOR U10828 ( .A(n10867), .B(n11013), .Z(n10860) );
  IV U10829 ( .A(n10866), .Z(n11013) );
  XNOR U10830 ( .A(n10863), .B(n11014), .Z(n10866) );
  XOR U10831 ( .A(n11015), .B(n11016), .Z(n10863) );
  ANDN U10832 ( .A(n11017), .B(n11018), .Z(n11016) );
  XNOR U10833 ( .A(n11015), .B(n11019), .Z(n11017) );
  XOR U10834 ( .A(n10874), .B(n11020), .Z(n10867) );
  IV U10835 ( .A(n10873), .Z(n11020) );
  XNOR U10836 ( .A(n10870), .B(n11021), .Z(n10873) );
  XOR U10837 ( .A(n11022), .B(n11023), .Z(n10870) );
  ANDN U10838 ( .A(n11024), .B(n11025), .Z(n11023) );
  XNOR U10839 ( .A(n11022), .B(n11026), .Z(n11024) );
  XOR U10840 ( .A(n10881), .B(n11027), .Z(n10874) );
  IV U10841 ( .A(n10880), .Z(n11027) );
  XNOR U10842 ( .A(n10877), .B(n11028), .Z(n10880) );
  XOR U10843 ( .A(n11029), .B(n11030), .Z(n10877) );
  ANDN U10844 ( .A(n11031), .B(n11032), .Z(n11030) );
  XNOR U10845 ( .A(n11029), .B(n11033), .Z(n11031) );
  XOR U10846 ( .A(n10888), .B(n11034), .Z(n10881) );
  IV U10847 ( .A(n10887), .Z(n11034) );
  XNOR U10848 ( .A(n10884), .B(n11035), .Z(n10887) );
  XOR U10849 ( .A(n11036), .B(n11037), .Z(n10884) );
  ANDN U10850 ( .A(n11038), .B(n11039), .Z(n11037) );
  XNOR U10851 ( .A(n11036), .B(n11040), .Z(n11038) );
  XOR U10852 ( .A(n10895), .B(n11041), .Z(n10888) );
  IV U10853 ( .A(n10894), .Z(n11041) );
  XNOR U10854 ( .A(n10891), .B(n11042), .Z(n10894) );
  XOR U10855 ( .A(n11043), .B(n11044), .Z(n10891) );
  ANDN U10856 ( .A(n11045), .B(n11046), .Z(n11044) );
  XNOR U10857 ( .A(n11043), .B(n11047), .Z(n11045) );
  XOR U10858 ( .A(n10901), .B(n11048), .Z(n10895) );
  IV U10859 ( .A(n10900), .Z(n11048) );
  XNOR U10860 ( .A(n10897), .B(n11049), .Z(n10900) );
  XOR U10861 ( .A(n11050), .B(n11051), .Z(n10897) );
  ANDN U10862 ( .A(n11052), .B(n11053), .Z(n11051) );
  XNOR U10863 ( .A(n11050), .B(n11054), .Z(n11052) );
  XOR U10864 ( .A(n10907), .B(n11055), .Z(n10901) );
  IV U10865 ( .A(n10906), .Z(n11055) );
  XNOR U10866 ( .A(n10903), .B(n11042), .Z(n10906) );
  AND U10867 ( .A(n11341), .B(n10731), .Z(n11042) );
  XOR U10868 ( .A(n11056), .B(n11057), .Z(n10903) );
  ANDN U10869 ( .A(n11058), .B(n11059), .Z(n11057) );
  XNOR U10870 ( .A(n11056), .B(n11060), .Z(n11058) );
  XOR U10871 ( .A(n10913), .B(n11061), .Z(n10907) );
  IV U10872 ( .A(n10912), .Z(n11061) );
  XNOR U10873 ( .A(n10909), .B(n11035), .Z(n10912) );
  AND U10874 ( .A(n11607), .B(n10387), .Z(n11035) );
  XOR U10875 ( .A(n11062), .B(n11063), .Z(n10909) );
  ANDN U10876 ( .A(n11064), .B(n11065), .Z(n11063) );
  XNOR U10877 ( .A(n11062), .B(n11066), .Z(n11064) );
  XOR U10878 ( .A(n10919), .B(n11067), .Z(n10913) );
  IV U10879 ( .A(n10918), .Z(n11067) );
  XNOR U10880 ( .A(n10915), .B(n11028), .Z(n10918) );
  AND U10881 ( .A(n11869), .B(n10017), .Z(n11028) );
  XOR U10882 ( .A(n11068), .B(n11069), .Z(n10915) );
  ANDN U10883 ( .A(n11070), .B(n11071), .Z(n11069) );
  XNOR U10884 ( .A(n11068), .B(n11072), .Z(n11070) );
  XOR U10885 ( .A(n10925), .B(n11073), .Z(n10919) );
  IV U10886 ( .A(n10924), .Z(n11073) );
  XNOR U10887 ( .A(n10921), .B(n11021), .Z(n10924) );
  AND U10888 ( .A(n12128), .B(n9621), .Z(n11021) );
  XOR U10889 ( .A(n11074), .B(n11075), .Z(n10921) );
  ANDN U10890 ( .A(n11076), .B(n11077), .Z(n11075) );
  XNOR U10891 ( .A(n11074), .B(n11078), .Z(n11076) );
  XOR U10892 ( .A(n10931), .B(n11079), .Z(n10925) );
  IV U10893 ( .A(n10930), .Z(n11079) );
  XNOR U10894 ( .A(n10927), .B(n11014), .Z(n10930) );
  AND U10895 ( .A(n12387), .B(n9198), .Z(n11014) );
  XOR U10896 ( .A(n11080), .B(n11081), .Z(n10927) );
  ANDN U10897 ( .A(n11082), .B(n11083), .Z(n11081) );
  XNOR U10898 ( .A(n11080), .B(n11084), .Z(n11082) );
  XOR U10899 ( .A(n10937), .B(n11085), .Z(n10931) );
  IV U10900 ( .A(n10936), .Z(n11085) );
  XNOR U10901 ( .A(n10933), .B(n11007), .Z(n10936) );
  AND U10902 ( .A(n12644), .B(n8748), .Z(n11007) );
  XOR U10903 ( .A(n11086), .B(n11087), .Z(n10933) );
  ANDN U10904 ( .A(n11088), .B(n11089), .Z(n11087) );
  XNOR U10905 ( .A(n11086), .B(n11090), .Z(n11088) );
  XOR U10906 ( .A(n10943), .B(n11091), .Z(n10937) );
  IV U10907 ( .A(n10942), .Z(n11091) );
  XNOR U10908 ( .A(n10939), .B(n11000), .Z(n10942) );
  AND U10909 ( .A(n12880), .B(n8272), .Z(n11000) );
  XOR U10910 ( .A(n11092), .B(n11093), .Z(n10939) );
  ANDN U10911 ( .A(n11094), .B(n11095), .Z(n11093) );
  XNOR U10912 ( .A(n11092), .B(n11096), .Z(n11094) );
  XOR U10913 ( .A(n10949), .B(n11097), .Z(n10943) );
  IV U10914 ( .A(n10948), .Z(n11097) );
  XNOR U10915 ( .A(n10945), .B(n10993), .Z(n10948) );
  AND U10916 ( .A(n13070), .B(n7770), .Z(n10993) );
  XOR U10917 ( .A(n11098), .B(n11099), .Z(n10945) );
  ANDN U10918 ( .A(n11100), .B(n11101), .Z(n11099) );
  XNOR U10919 ( .A(n11098), .B(n11102), .Z(n11100) );
  XOR U10920 ( .A(n10955), .B(n11103), .Z(n10949) );
  IV U10921 ( .A(n10954), .Z(n11103) );
  XNOR U10922 ( .A(n10951), .B(n10986), .Z(n10954) );
  AND U10923 ( .A(n13207), .B(n7241), .Z(n10986) );
  XOR U10924 ( .A(n11104), .B(n11105), .Z(n10951) );
  ANDN U10925 ( .A(n11106), .B(n11107), .Z(n11105) );
  XNOR U10926 ( .A(n11104), .B(n11108), .Z(n11106) );
  XNOR U10927 ( .A(n10960), .B(n10824), .Z(n10955) );
  XNOR U10928 ( .A(n10957), .B(n11109), .Z(n10960) );
  AND U10929 ( .A(n6527), .B(n6688), .Z(n11109) );
  XOR U10930 ( .A(n11110), .B(n11111), .Z(n10957) );
  ANDN U10931 ( .A(n11112), .B(n11113), .Z(n11111) );
  XNOR U10932 ( .A(n10983), .B(n11110), .Z(n11112) );
  XOR U10933 ( .A(n11114), .B(n10824), .Z(n10980) );
  NANDN U10934 ( .B(n6808), .A(n6118), .Z(n10824) );
  XOR U10935 ( .A(n11115), .B(n11116), .Z(n6118) );
  AND U10936 ( .A(n6809), .B(n11117), .Z(n11116) );
  XNOR U10937 ( .A(n11115), .B(n10967), .Z(n11117) );
  XOR U10938 ( .A(n10965), .B(n11115), .Z(n10967) );
  XOR U10939 ( .A(n11118), .B(n11119), .Z(n10965) );
  ANDN U10940 ( .A(n11118), .B(n11120), .Z(n11119) );
  XOR U10941 ( .A(n11121), .B(n7368), .Z(n11115) );
  IV U10942 ( .A(n10969), .Z(n11114) );
  XOR U10943 ( .A(n11122), .B(n11123), .Z(n10969) );
  AND U10944 ( .A(n11124), .B(n11125), .Z(n11123) );
  XNOR U10945 ( .A(n11126), .B(n11122), .Z(n11125) );
  XNOR U10946 ( .A(n10973), .B(n10976), .Z(n10979) );
  XOR U10947 ( .A(n11127), .B(n11128), .Z(n10973) );
  XOR U10948 ( .A(n11129), .B(n11130), .Z(n10976) );
  AND U10949 ( .A(n11129), .B(n11131), .Z(n11130) );
  XOR U10950 ( .A(n11132), .B(n11124), .Z(n11131) );
  XOR U10951 ( .A(n11133), .B(n10984), .Z(n11124) );
  XOR U10952 ( .A(n10991), .B(n11134), .Z(n10984) );
  IV U10953 ( .A(n10989), .Z(n11134) );
  XNOR U10954 ( .A(n11135), .B(n10988), .Z(n10989) );
  OR U10955 ( .A(n11136), .B(n11137), .Z(n10988) );
  NANDN U10956 ( .B(n6541), .A(n7241), .Z(n11135) );
  XOR U10957 ( .A(n10998), .B(n11138), .Z(n10991) );
  IV U10958 ( .A(n10997), .Z(n11138) );
  XNOR U10959 ( .A(n10994), .B(n11139), .Z(n10997) );
  XOR U10960 ( .A(n11140), .B(n11141), .Z(n10994) );
  NANDN U10961 ( .B(n11142), .A(n11143), .Z(n11140) );
  XOR U10962 ( .A(n11141), .B(n11144), .Z(n11143) );
  XOR U10963 ( .A(n11005), .B(n11145), .Z(n10998) );
  IV U10964 ( .A(n11004), .Z(n11145) );
  XNOR U10965 ( .A(n11001), .B(n11146), .Z(n11004) );
  XOR U10966 ( .A(n11147), .B(n11148), .Z(n11001) );
  ANDN U10967 ( .A(n11149), .B(n11150), .Z(n11148) );
  XNOR U10968 ( .A(n11147), .B(n11151), .Z(n11149) );
  XOR U10969 ( .A(n11012), .B(n11152), .Z(n11005) );
  IV U10970 ( .A(n11011), .Z(n11152) );
  XNOR U10971 ( .A(n11008), .B(n11153), .Z(n11011) );
  XOR U10972 ( .A(n11154), .B(n11155), .Z(n11008) );
  ANDN U10973 ( .A(n11156), .B(n11157), .Z(n11155) );
  XNOR U10974 ( .A(n11154), .B(n11158), .Z(n11156) );
  XOR U10975 ( .A(n11019), .B(n11159), .Z(n11012) );
  IV U10976 ( .A(n11018), .Z(n11159) );
  XNOR U10977 ( .A(n11015), .B(n11160), .Z(n11018) );
  XOR U10978 ( .A(n11161), .B(n11162), .Z(n11015) );
  ANDN U10979 ( .A(n11163), .B(n11164), .Z(n11162) );
  XNOR U10980 ( .A(n11161), .B(n11165), .Z(n11163) );
  XOR U10981 ( .A(n11026), .B(n11166), .Z(n11019) );
  IV U10982 ( .A(n11025), .Z(n11166) );
  XNOR U10983 ( .A(n11022), .B(n11167), .Z(n11025) );
  XOR U10984 ( .A(n11168), .B(n11169), .Z(n11022) );
  ANDN U10985 ( .A(n11170), .B(n11171), .Z(n11169) );
  XNOR U10986 ( .A(n11168), .B(n11172), .Z(n11170) );
  XOR U10987 ( .A(n11033), .B(n11173), .Z(n11026) );
  IV U10988 ( .A(n11032), .Z(n11173) );
  XNOR U10989 ( .A(n11029), .B(n11174), .Z(n11032) );
  XOR U10990 ( .A(n11175), .B(n11176), .Z(n11029) );
  ANDN U10991 ( .A(n11177), .B(n11178), .Z(n11176) );
  XNOR U10992 ( .A(n11175), .B(n11179), .Z(n11177) );
  XOR U10993 ( .A(n11040), .B(n11180), .Z(n11033) );
  IV U10994 ( .A(n11039), .Z(n11180) );
  XNOR U10995 ( .A(n11036), .B(n11181), .Z(n11039) );
  XOR U10996 ( .A(n11182), .B(n11183), .Z(n11036) );
  ANDN U10997 ( .A(n11184), .B(n11185), .Z(n11183) );
  XNOR U10998 ( .A(n11182), .B(n11186), .Z(n11184) );
  XOR U10999 ( .A(n11047), .B(n11187), .Z(n11040) );
  IV U11000 ( .A(n11046), .Z(n11187) );
  XNOR U11001 ( .A(n11043), .B(n11188), .Z(n11046) );
  XOR U11002 ( .A(n11189), .B(n11190), .Z(n11043) );
  ANDN U11003 ( .A(n11191), .B(n11192), .Z(n11190) );
  XNOR U11004 ( .A(n11189), .B(n11193), .Z(n11191) );
  XOR U11005 ( .A(n11054), .B(n11194), .Z(n11047) );
  IV U11006 ( .A(n11053), .Z(n11194) );
  XNOR U11007 ( .A(n11050), .B(n11195), .Z(n11053) );
  XOR U11008 ( .A(n11196), .B(n11197), .Z(n11050) );
  ANDN U11009 ( .A(n11198), .B(n11199), .Z(n11197) );
  XNOR U11010 ( .A(n11196), .B(n11200), .Z(n11198) );
  XOR U11011 ( .A(n11060), .B(n11201), .Z(n11054) );
  IV U11012 ( .A(n11059), .Z(n11201) );
  XNOR U11013 ( .A(n11056), .B(n11195), .Z(n11059) );
  AND U11014 ( .A(n11341), .B(n11049), .Z(n11195) );
  XOR U11015 ( .A(n11202), .B(n11203), .Z(n11056) );
  ANDN U11016 ( .A(n11204), .B(n11205), .Z(n11203) );
  XNOR U11017 ( .A(n11202), .B(n11206), .Z(n11204) );
  XOR U11018 ( .A(n11066), .B(n11207), .Z(n11060) );
  IV U11019 ( .A(n11065), .Z(n11207) );
  XNOR U11020 ( .A(n11062), .B(n11188), .Z(n11065) );
  AND U11021 ( .A(n11607), .B(n10731), .Z(n11188) );
  XOR U11022 ( .A(n11208), .B(n11209), .Z(n11062) );
  ANDN U11023 ( .A(n11210), .B(n11211), .Z(n11209) );
  XNOR U11024 ( .A(n11208), .B(n11212), .Z(n11210) );
  XOR U11025 ( .A(n11072), .B(n11213), .Z(n11066) );
  IV U11026 ( .A(n11071), .Z(n11213) );
  XNOR U11027 ( .A(n11068), .B(n11181), .Z(n11071) );
  AND U11028 ( .A(n11869), .B(n10387), .Z(n11181) );
  XOR U11029 ( .A(n11214), .B(n11215), .Z(n11068) );
  ANDN U11030 ( .A(n11216), .B(n11217), .Z(n11215) );
  XNOR U11031 ( .A(n11214), .B(n11218), .Z(n11216) );
  XOR U11032 ( .A(n11078), .B(n11219), .Z(n11072) );
  IV U11033 ( .A(n11077), .Z(n11219) );
  XNOR U11034 ( .A(n11074), .B(n11174), .Z(n11077) );
  AND U11035 ( .A(n12128), .B(n10017), .Z(n11174) );
  XOR U11036 ( .A(n11220), .B(n11221), .Z(n11074) );
  ANDN U11037 ( .A(n11222), .B(n11223), .Z(n11221) );
  XNOR U11038 ( .A(n11220), .B(n11224), .Z(n11222) );
  XOR U11039 ( .A(n11084), .B(n11225), .Z(n11078) );
  IV U11040 ( .A(n11083), .Z(n11225) );
  XNOR U11041 ( .A(n11080), .B(n11167), .Z(n11083) );
  AND U11042 ( .A(n12387), .B(n9621), .Z(n11167) );
  XOR U11043 ( .A(n11226), .B(n11227), .Z(n11080) );
  ANDN U11044 ( .A(n11228), .B(n11229), .Z(n11227) );
  XNOR U11045 ( .A(n11226), .B(n11230), .Z(n11228) );
  XOR U11046 ( .A(n11090), .B(n11231), .Z(n11084) );
  IV U11047 ( .A(n11089), .Z(n11231) );
  XNOR U11048 ( .A(n11086), .B(n11160), .Z(n11089) );
  AND U11049 ( .A(n12644), .B(n9198), .Z(n11160) );
  XOR U11050 ( .A(n11232), .B(n11233), .Z(n11086) );
  ANDN U11051 ( .A(n11234), .B(n11235), .Z(n11233) );
  XNOR U11052 ( .A(n11232), .B(n11236), .Z(n11234) );
  XOR U11053 ( .A(n11096), .B(n11237), .Z(n11090) );
  IV U11054 ( .A(n11095), .Z(n11237) );
  XNOR U11055 ( .A(n11092), .B(n11153), .Z(n11095) );
  AND U11056 ( .A(n12880), .B(n8748), .Z(n11153) );
  XOR U11057 ( .A(n11238), .B(n11239), .Z(n11092) );
  ANDN U11058 ( .A(n11240), .B(n11241), .Z(n11239) );
  XNOR U11059 ( .A(n11238), .B(n11242), .Z(n11240) );
  XOR U11060 ( .A(n11102), .B(n11243), .Z(n11096) );
  IV U11061 ( .A(n11101), .Z(n11243) );
  XNOR U11062 ( .A(n11098), .B(n11146), .Z(n11101) );
  AND U11063 ( .A(n13070), .B(n8272), .Z(n11146) );
  XOR U11064 ( .A(n11244), .B(n11245), .Z(n11098) );
  ANDN U11065 ( .A(n11246), .B(n11247), .Z(n11245) );
  XNOR U11066 ( .A(n11244), .B(n11248), .Z(n11246) );
  XOR U11067 ( .A(n11108), .B(n11249), .Z(n11102) );
  IV U11068 ( .A(n11107), .Z(n11249) );
  XNOR U11069 ( .A(n11104), .B(n11139), .Z(n11107) );
  AND U11070 ( .A(n13207), .B(n7770), .Z(n11139) );
  XOR U11071 ( .A(n11250), .B(n11251), .Z(n11104) );
  ANDN U11072 ( .A(n11252), .B(n11253), .Z(n11251) );
  XNOR U11073 ( .A(n11250), .B(n11254), .Z(n11252) );
  XNOR U11074 ( .A(n11113), .B(n10983), .Z(n11108) );
  XNOR U11075 ( .A(n11110), .B(n11255), .Z(n11113) );
  AND U11076 ( .A(n6527), .B(n7241), .Z(n11255) );
  XOR U11077 ( .A(n11256), .B(n11257), .Z(n11110) );
  ANDN U11078 ( .A(n11258), .B(n11259), .Z(n11257) );
  XNOR U11079 ( .A(n11136), .B(n11256), .Z(n11258) );
  XOR U11080 ( .A(n11260), .B(n10983), .Z(n11133) );
  NANDN U11081 ( .B(n6808), .A(n6688), .Z(n10983) );
  XOR U11082 ( .A(n11261), .B(n11262), .Z(n6688) );
  AND U11083 ( .A(n6809), .B(n11263), .Z(n11262) );
  XNOR U11084 ( .A(n11261), .B(n11120), .Z(n11263) );
  XOR U11085 ( .A(n11118), .B(n11261), .Z(n11120) );
  XOR U11086 ( .A(n11264), .B(n11265), .Z(n11118) );
  ANDN U11087 ( .A(n11264), .B(n11266), .Z(n11265) );
  XOR U11088 ( .A(n11267), .B(n7368), .Z(n11261) );
  IV U11089 ( .A(n11122), .Z(n11260) );
  XOR U11090 ( .A(n11268), .B(n11269), .Z(n11122) );
  AND U11091 ( .A(n11270), .B(n11271), .Z(n11269) );
  XNOR U11092 ( .A(n11272), .B(n11268), .Z(n11271) );
  XNOR U11093 ( .A(n11126), .B(n11129), .Z(n11132) );
  XOR U11094 ( .A(n11273), .B(n11274), .Z(n11126) );
  XOR U11095 ( .A(n11275), .B(n11276), .Z(n11129) );
  AND U11096 ( .A(n11275), .B(n11277), .Z(n11276) );
  XOR U11097 ( .A(n11278), .B(n11270), .Z(n11277) );
  XOR U11098 ( .A(n11279), .B(n11137), .Z(n11270) );
  XOR U11099 ( .A(n11144), .B(n11280), .Z(n11137) );
  IV U11100 ( .A(n11142), .Z(n11280) );
  XNOR U11101 ( .A(n11281), .B(n11141), .Z(n11142) );
  OR U11102 ( .A(n11282), .B(n11283), .Z(n11141) );
  NANDN U11103 ( .B(n6541), .A(n7770), .Z(n11281) );
  XOR U11104 ( .A(n11151), .B(n11284), .Z(n11144) );
  IV U11105 ( .A(n11150), .Z(n11284) );
  XNOR U11106 ( .A(n11147), .B(n11285), .Z(n11150) );
  XOR U11107 ( .A(n11286), .B(n11287), .Z(n11147) );
  NANDN U11108 ( .B(n11288), .A(n11289), .Z(n11286) );
  XOR U11109 ( .A(n11287), .B(n11290), .Z(n11289) );
  XOR U11110 ( .A(n11158), .B(n11291), .Z(n11151) );
  IV U11111 ( .A(n11157), .Z(n11291) );
  XNOR U11112 ( .A(n11154), .B(n11292), .Z(n11157) );
  XOR U11113 ( .A(n11293), .B(n11294), .Z(n11154) );
  ANDN U11114 ( .A(n11295), .B(n11296), .Z(n11294) );
  XNOR U11115 ( .A(n11293), .B(n11297), .Z(n11295) );
  XOR U11116 ( .A(n11165), .B(n11298), .Z(n11158) );
  IV U11117 ( .A(n11164), .Z(n11298) );
  XNOR U11118 ( .A(n11161), .B(n11299), .Z(n11164) );
  XOR U11119 ( .A(n11300), .B(n11301), .Z(n11161) );
  ANDN U11120 ( .A(n11302), .B(n11303), .Z(n11301) );
  XNOR U11121 ( .A(n11300), .B(n11304), .Z(n11302) );
  XOR U11122 ( .A(n11172), .B(n11305), .Z(n11165) );
  IV U11123 ( .A(n11171), .Z(n11305) );
  XNOR U11124 ( .A(n11168), .B(n11306), .Z(n11171) );
  XOR U11125 ( .A(n11307), .B(n11308), .Z(n11168) );
  ANDN U11126 ( .A(n11309), .B(n11310), .Z(n11308) );
  XNOR U11127 ( .A(n11307), .B(n11311), .Z(n11309) );
  XOR U11128 ( .A(n11179), .B(n11312), .Z(n11172) );
  IV U11129 ( .A(n11178), .Z(n11312) );
  XNOR U11130 ( .A(n11175), .B(n11313), .Z(n11178) );
  XOR U11131 ( .A(n11314), .B(n11315), .Z(n11175) );
  ANDN U11132 ( .A(n11316), .B(n11317), .Z(n11315) );
  XNOR U11133 ( .A(n11314), .B(n11318), .Z(n11316) );
  XOR U11134 ( .A(n11186), .B(n11319), .Z(n11179) );
  IV U11135 ( .A(n11185), .Z(n11319) );
  XNOR U11136 ( .A(n11182), .B(n11320), .Z(n11185) );
  XOR U11137 ( .A(n11321), .B(n11322), .Z(n11182) );
  ANDN U11138 ( .A(n11323), .B(n11324), .Z(n11322) );
  XNOR U11139 ( .A(n11321), .B(n11325), .Z(n11323) );
  XOR U11140 ( .A(n11193), .B(n11326), .Z(n11186) );
  IV U11141 ( .A(n11192), .Z(n11326) );
  XNOR U11142 ( .A(n11189), .B(n11327), .Z(n11192) );
  XOR U11143 ( .A(n11328), .B(n11329), .Z(n11189) );
  ANDN U11144 ( .A(n11330), .B(n11331), .Z(n11329) );
  XNOR U11145 ( .A(n11328), .B(n11332), .Z(n11330) );
  XOR U11146 ( .A(n11200), .B(n11333), .Z(n11193) );
  IV U11147 ( .A(n11199), .Z(n11333) );
  XNOR U11148 ( .A(n11196), .B(n11334), .Z(n11199) );
  XOR U11149 ( .A(n11335), .B(n11336), .Z(n11196) );
  ANDN U11150 ( .A(n11337), .B(n11338), .Z(n11336) );
  XNOR U11151 ( .A(n11335), .B(n11339), .Z(n11337) );
  XOR U11152 ( .A(n11206), .B(n11340), .Z(n11200) );
  IV U11153 ( .A(n11205), .Z(n11340) );
  XNOR U11154 ( .A(n11202), .B(n11341), .Z(n11205) );
  XOR U11155 ( .A(n11342), .B(n11343), .Z(n11202) );
  ANDN U11156 ( .A(n11344), .B(n11345), .Z(n11343) );
  XNOR U11157 ( .A(n11342), .B(n11346), .Z(n11344) );
  XOR U11158 ( .A(n11212), .B(n11347), .Z(n11206) );
  IV U11159 ( .A(n11211), .Z(n11347) );
  XNOR U11160 ( .A(n11208), .B(n11334), .Z(n11211) );
  AND U11161 ( .A(n11607), .B(n11049), .Z(n11334) );
  XOR U11162 ( .A(n11348), .B(n11349), .Z(n11208) );
  ANDN U11163 ( .A(n11350), .B(n11351), .Z(n11349) );
  XNOR U11164 ( .A(n11348), .B(n11352), .Z(n11350) );
  XOR U11165 ( .A(n11218), .B(n11353), .Z(n11212) );
  IV U11166 ( .A(n11217), .Z(n11353) );
  XNOR U11167 ( .A(n11214), .B(n11327), .Z(n11217) );
  AND U11168 ( .A(n11869), .B(n10731), .Z(n11327) );
  XOR U11169 ( .A(n11354), .B(n11355), .Z(n11214) );
  ANDN U11170 ( .A(n11356), .B(n11357), .Z(n11355) );
  XNOR U11171 ( .A(n11354), .B(n11358), .Z(n11356) );
  XOR U11172 ( .A(n11224), .B(n11359), .Z(n11218) );
  IV U11173 ( .A(n11223), .Z(n11359) );
  XNOR U11174 ( .A(n11220), .B(n11320), .Z(n11223) );
  AND U11175 ( .A(n12128), .B(n10387), .Z(n11320) );
  XOR U11176 ( .A(n11360), .B(n11361), .Z(n11220) );
  ANDN U11177 ( .A(n11362), .B(n11363), .Z(n11361) );
  XNOR U11178 ( .A(n11360), .B(n11364), .Z(n11362) );
  XOR U11179 ( .A(n11230), .B(n11365), .Z(n11224) );
  IV U11180 ( .A(n11229), .Z(n11365) );
  XNOR U11181 ( .A(n11226), .B(n11313), .Z(n11229) );
  AND U11182 ( .A(n12387), .B(n10017), .Z(n11313) );
  XOR U11183 ( .A(n11366), .B(n11367), .Z(n11226) );
  ANDN U11184 ( .A(n11368), .B(n11369), .Z(n11367) );
  XNOR U11185 ( .A(n11366), .B(n11370), .Z(n11368) );
  XOR U11186 ( .A(n11236), .B(n11371), .Z(n11230) );
  IV U11187 ( .A(n11235), .Z(n11371) );
  XNOR U11188 ( .A(n11232), .B(n11306), .Z(n11235) );
  AND U11189 ( .A(n12644), .B(n9621), .Z(n11306) );
  XOR U11190 ( .A(n11372), .B(n11373), .Z(n11232) );
  ANDN U11191 ( .A(n11374), .B(n11375), .Z(n11373) );
  XNOR U11192 ( .A(n11372), .B(n11376), .Z(n11374) );
  XOR U11193 ( .A(n11242), .B(n11377), .Z(n11236) );
  IV U11194 ( .A(n11241), .Z(n11377) );
  XNOR U11195 ( .A(n11238), .B(n11299), .Z(n11241) );
  AND U11196 ( .A(n12880), .B(n9198), .Z(n11299) );
  XOR U11197 ( .A(n11378), .B(n11379), .Z(n11238) );
  ANDN U11198 ( .A(n11380), .B(n11381), .Z(n11379) );
  XNOR U11199 ( .A(n11378), .B(n11382), .Z(n11380) );
  XOR U11200 ( .A(n11248), .B(n11383), .Z(n11242) );
  IV U11201 ( .A(n11247), .Z(n11383) );
  XNOR U11202 ( .A(n11244), .B(n11292), .Z(n11247) );
  AND U11203 ( .A(n13070), .B(n8748), .Z(n11292) );
  XOR U11204 ( .A(n11384), .B(n11385), .Z(n11244) );
  ANDN U11205 ( .A(n11386), .B(n11387), .Z(n11385) );
  XNOR U11206 ( .A(n11384), .B(n11388), .Z(n11386) );
  XOR U11207 ( .A(n11254), .B(n11389), .Z(n11248) );
  IV U11208 ( .A(n11253), .Z(n11389) );
  XNOR U11209 ( .A(n11250), .B(n11285), .Z(n11253) );
  AND U11210 ( .A(n13207), .B(n8272), .Z(n11285) );
  XOR U11211 ( .A(n11390), .B(n11391), .Z(n11250) );
  ANDN U11212 ( .A(n11392), .B(n11393), .Z(n11391) );
  XNOR U11213 ( .A(n11390), .B(n11394), .Z(n11392) );
  XNOR U11214 ( .A(n11259), .B(n11136), .Z(n11254) );
  XNOR U11215 ( .A(n11256), .B(n11395), .Z(n11259) );
  AND U11216 ( .A(n6527), .B(n7770), .Z(n11395) );
  XOR U11217 ( .A(n11396), .B(n11397), .Z(n11256) );
  ANDN U11218 ( .A(n11398), .B(n11399), .Z(n11397) );
  XNOR U11219 ( .A(n11282), .B(n11396), .Z(n11398) );
  XOR U11220 ( .A(n11400), .B(n11136), .Z(n11279) );
  NANDN U11221 ( .B(n6808), .A(n7241), .Z(n11136) );
  XOR U11222 ( .A(n11401), .B(n11402), .Z(n7241) );
  AND U11223 ( .A(n6809), .B(n11403), .Z(n11402) );
  XNOR U11224 ( .A(n11401), .B(n11266), .Z(n11403) );
  XOR U11225 ( .A(n11264), .B(n11401), .Z(n11266) );
  XOR U11226 ( .A(n11404), .B(n11405), .Z(n11264) );
  ANDN U11227 ( .A(n11404), .B(n11406), .Z(n11405) );
  XOR U11228 ( .A(n11407), .B(n7368), .Z(n11401) );
  IV U11229 ( .A(n11268), .Z(n11400) );
  XOR U11230 ( .A(n11408), .B(n11409), .Z(n11268) );
  AND U11231 ( .A(n11410), .B(n11411), .Z(n11409) );
  XNOR U11232 ( .A(n11412), .B(n11408), .Z(n11411) );
  XNOR U11233 ( .A(n11272), .B(n11275), .Z(n11278) );
  XOR U11234 ( .A(n11413), .B(n11414), .Z(n11272) );
  XOR U11235 ( .A(n11415), .B(n11416), .Z(n11275) );
  AND U11236 ( .A(n11415), .B(n11417), .Z(n11416) );
  XOR U11237 ( .A(n11418), .B(n11410), .Z(n11417) );
  XOR U11238 ( .A(n11419), .B(n11283), .Z(n11410) );
  XOR U11239 ( .A(n11290), .B(n11420), .Z(n11283) );
  IV U11240 ( .A(n11288), .Z(n11420) );
  XNOR U11241 ( .A(n11421), .B(n11287), .Z(n11288) );
  OR U11242 ( .A(n11422), .B(n11423), .Z(n11287) );
  NANDN U11243 ( .B(n6541), .A(n8272), .Z(n11421) );
  XOR U11244 ( .A(n11297), .B(n11424), .Z(n11290) );
  IV U11245 ( .A(n11296), .Z(n11424) );
  XNOR U11246 ( .A(n11293), .B(n11425), .Z(n11296) );
  XOR U11247 ( .A(n11426), .B(n11427), .Z(n11293) );
  NANDN U11248 ( .B(n11428), .A(n11429), .Z(n11426) );
  XOR U11249 ( .A(n11427), .B(n11430), .Z(n11429) );
  XOR U11250 ( .A(n11304), .B(n11431), .Z(n11297) );
  IV U11251 ( .A(n11303), .Z(n11431) );
  XNOR U11252 ( .A(n11300), .B(n11432), .Z(n11303) );
  XOR U11253 ( .A(n11433), .B(n11434), .Z(n11300) );
  ANDN U11254 ( .A(n11435), .B(n11436), .Z(n11434) );
  XNOR U11255 ( .A(n11433), .B(n11437), .Z(n11435) );
  XOR U11256 ( .A(n11311), .B(n11438), .Z(n11304) );
  IV U11257 ( .A(n11310), .Z(n11438) );
  XNOR U11258 ( .A(n11307), .B(n11439), .Z(n11310) );
  XOR U11259 ( .A(n11440), .B(n11441), .Z(n11307) );
  ANDN U11260 ( .A(n11442), .B(n11443), .Z(n11441) );
  XNOR U11261 ( .A(n11440), .B(n11444), .Z(n11442) );
  XOR U11262 ( .A(n11318), .B(n11445), .Z(n11311) );
  IV U11263 ( .A(n11317), .Z(n11445) );
  XNOR U11264 ( .A(n11314), .B(n11446), .Z(n11317) );
  XOR U11265 ( .A(n11447), .B(n11448), .Z(n11314) );
  ANDN U11266 ( .A(n11449), .B(n11450), .Z(n11448) );
  XNOR U11267 ( .A(n11447), .B(n11451), .Z(n11449) );
  XOR U11268 ( .A(n11325), .B(n11452), .Z(n11318) );
  IV U11269 ( .A(n11324), .Z(n11452) );
  XNOR U11270 ( .A(n11321), .B(n11453), .Z(n11324) );
  XOR U11271 ( .A(n11454), .B(n11455), .Z(n11321) );
  ANDN U11272 ( .A(n11456), .B(n11457), .Z(n11455) );
  XNOR U11273 ( .A(n11454), .B(n11458), .Z(n11456) );
  XOR U11274 ( .A(n11332), .B(n11459), .Z(n11325) );
  IV U11275 ( .A(n11331), .Z(n11459) );
  XNOR U11276 ( .A(n11328), .B(n11460), .Z(n11331) );
  XOR U11277 ( .A(n11461), .B(n11462), .Z(n11328) );
  ANDN U11278 ( .A(n11463), .B(n11464), .Z(n11462) );
  XNOR U11279 ( .A(n11461), .B(n11465), .Z(n11463) );
  XOR U11280 ( .A(n11339), .B(n11466), .Z(n11332) );
  IV U11281 ( .A(n11338), .Z(n11466) );
  XNOR U11282 ( .A(n11335), .B(n11467), .Z(n11338) );
  XOR U11283 ( .A(n11468), .B(n11469), .Z(n11335) );
  ANDN U11284 ( .A(n11470), .B(n11471), .Z(n11469) );
  XNOR U11285 ( .A(n11468), .B(n11472), .Z(n11470) );
  XOR U11286 ( .A(n11346), .B(n11473), .Z(n11339) );
  IV U11287 ( .A(n11345), .Z(n11473) );
  XNOR U11288 ( .A(n11342), .B(n11474), .Z(n11345) );
  XOR U11289 ( .A(n11475), .B(n11476), .Z(n11342) );
  ANDN U11290 ( .A(n11477), .B(n11478), .Z(n11476) );
  XNOR U11291 ( .A(n11475), .B(n11479), .Z(n11477) );
  XOR U11292 ( .A(n11352), .B(n11480), .Z(n11346) );
  IV U11293 ( .A(n11351), .Z(n11480) );
  XNOR U11294 ( .A(n11348), .B(n11474), .Z(n11351) );
  AND U11295 ( .A(n11607), .B(n11341), .Z(n11474) );
  XOR U11296 ( .A(n11481), .B(n11482), .Z(n11348) );
  ANDN U11297 ( .A(n11483), .B(n11484), .Z(n11482) );
  XNOR U11298 ( .A(n11481), .B(n11485), .Z(n11483) );
  XOR U11299 ( .A(n11358), .B(n11486), .Z(n11352) );
  IV U11300 ( .A(n11357), .Z(n11486) );
  XNOR U11301 ( .A(n11354), .B(n11467), .Z(n11357) );
  AND U11302 ( .A(n11869), .B(n11049), .Z(n11467) );
  XOR U11303 ( .A(n11487), .B(n11488), .Z(n11354) );
  ANDN U11304 ( .A(n11489), .B(n11490), .Z(n11488) );
  XNOR U11305 ( .A(n11487), .B(n11491), .Z(n11489) );
  XOR U11306 ( .A(n11364), .B(n11492), .Z(n11358) );
  IV U11307 ( .A(n11363), .Z(n11492) );
  XNOR U11308 ( .A(n11360), .B(n11460), .Z(n11363) );
  AND U11309 ( .A(n12128), .B(n10731), .Z(n11460) );
  XOR U11310 ( .A(n11493), .B(n11494), .Z(n11360) );
  ANDN U11311 ( .A(n11495), .B(n11496), .Z(n11494) );
  XNOR U11312 ( .A(n11493), .B(n11497), .Z(n11495) );
  XOR U11313 ( .A(n11370), .B(n11498), .Z(n11364) );
  IV U11314 ( .A(n11369), .Z(n11498) );
  XNOR U11315 ( .A(n11366), .B(n11453), .Z(n11369) );
  AND U11316 ( .A(n12387), .B(n10387), .Z(n11453) );
  XOR U11317 ( .A(n11499), .B(n11500), .Z(n11366) );
  ANDN U11318 ( .A(n11501), .B(n11502), .Z(n11500) );
  XNOR U11319 ( .A(n11499), .B(n11503), .Z(n11501) );
  XOR U11320 ( .A(n11376), .B(n11504), .Z(n11370) );
  IV U11321 ( .A(n11375), .Z(n11504) );
  XNOR U11322 ( .A(n11372), .B(n11446), .Z(n11375) );
  AND U11323 ( .A(n12644), .B(n10017), .Z(n11446) );
  XOR U11324 ( .A(n11505), .B(n11506), .Z(n11372) );
  ANDN U11325 ( .A(n11507), .B(n11508), .Z(n11506) );
  XNOR U11326 ( .A(n11505), .B(n11509), .Z(n11507) );
  XOR U11327 ( .A(n11382), .B(n11510), .Z(n11376) );
  IV U11328 ( .A(n11381), .Z(n11510) );
  XNOR U11329 ( .A(n11378), .B(n11439), .Z(n11381) );
  AND U11330 ( .A(n12880), .B(n9621), .Z(n11439) );
  XOR U11331 ( .A(n11511), .B(n11512), .Z(n11378) );
  ANDN U11332 ( .A(n11513), .B(n11514), .Z(n11512) );
  XNOR U11333 ( .A(n11511), .B(n11515), .Z(n11513) );
  XOR U11334 ( .A(n11388), .B(n11516), .Z(n11382) );
  IV U11335 ( .A(n11387), .Z(n11516) );
  XNOR U11336 ( .A(n11384), .B(n11432), .Z(n11387) );
  AND U11337 ( .A(n13070), .B(n9198), .Z(n11432) );
  XOR U11338 ( .A(n11517), .B(n11518), .Z(n11384) );
  ANDN U11339 ( .A(n11519), .B(n11520), .Z(n11518) );
  XNOR U11340 ( .A(n11517), .B(n11521), .Z(n11519) );
  XOR U11341 ( .A(n11394), .B(n11522), .Z(n11388) );
  IV U11342 ( .A(n11393), .Z(n11522) );
  XNOR U11343 ( .A(n11390), .B(n11425), .Z(n11393) );
  AND U11344 ( .A(n13207), .B(n8748), .Z(n11425) );
  XOR U11345 ( .A(n11523), .B(n11524), .Z(n11390) );
  ANDN U11346 ( .A(n11525), .B(n11526), .Z(n11524) );
  XNOR U11347 ( .A(n11523), .B(n11527), .Z(n11525) );
  XNOR U11348 ( .A(n11399), .B(n11282), .Z(n11394) );
  XNOR U11349 ( .A(n11396), .B(n11528), .Z(n11399) );
  AND U11350 ( .A(n6527), .B(n8272), .Z(n11528) );
  XOR U11351 ( .A(n11529), .B(n11530), .Z(n11396) );
  ANDN U11352 ( .A(n11531), .B(n11532), .Z(n11530) );
  XNOR U11353 ( .A(n11422), .B(n11529), .Z(n11531) );
  XOR U11354 ( .A(n11533), .B(n11282), .Z(n11419) );
  NANDN U11355 ( .B(n6808), .A(n7770), .Z(n11282) );
  XOR U11356 ( .A(n11534), .B(n11535), .Z(n7770) );
  AND U11357 ( .A(n6809), .B(n11536), .Z(n11535) );
  XNOR U11358 ( .A(n11534), .B(n11406), .Z(n11536) );
  XOR U11359 ( .A(n11404), .B(n11534), .Z(n11406) );
  XOR U11360 ( .A(n11537), .B(n11538), .Z(n11404) );
  ANDN U11361 ( .A(n11537), .B(n11539), .Z(n11538) );
  XOR U11362 ( .A(n11540), .B(n7368), .Z(n11534) );
  IV U11363 ( .A(n11408), .Z(n11533) );
  XOR U11364 ( .A(n11541), .B(n11542), .Z(n11408) );
  AND U11365 ( .A(n11543), .B(n11544), .Z(n11542) );
  XNOR U11366 ( .A(n11545), .B(n11541), .Z(n11544) );
  XNOR U11367 ( .A(n11412), .B(n11415), .Z(n11418) );
  XOR U11368 ( .A(n11546), .B(n11547), .Z(n11412) );
  XOR U11369 ( .A(n11548), .B(n11549), .Z(n11415) );
  AND U11370 ( .A(n11548), .B(n11550), .Z(n11549) );
  XOR U11371 ( .A(n11551), .B(n11543), .Z(n11550) );
  XOR U11372 ( .A(n11552), .B(n11423), .Z(n11543) );
  XOR U11373 ( .A(n11430), .B(n11553), .Z(n11423) );
  IV U11374 ( .A(n11428), .Z(n11553) );
  XNOR U11375 ( .A(n11554), .B(n11427), .Z(n11428) );
  OR U11376 ( .A(n11555), .B(n11556), .Z(n11427) );
  NANDN U11377 ( .B(n6541), .A(n8748), .Z(n11554) );
  XOR U11378 ( .A(n11437), .B(n11557), .Z(n11430) );
  IV U11379 ( .A(n11436), .Z(n11557) );
  XNOR U11380 ( .A(n11433), .B(n11558), .Z(n11436) );
  XOR U11381 ( .A(n11559), .B(n11560), .Z(n11433) );
  NANDN U11382 ( .B(n11561), .A(n11562), .Z(n11559) );
  XOR U11383 ( .A(n11560), .B(n11563), .Z(n11562) );
  XOR U11384 ( .A(n11444), .B(n11564), .Z(n11437) );
  IV U11385 ( .A(n11443), .Z(n11564) );
  XNOR U11386 ( .A(n11440), .B(n11565), .Z(n11443) );
  XOR U11387 ( .A(n11566), .B(n11567), .Z(n11440) );
  ANDN U11388 ( .A(n11568), .B(n11569), .Z(n11567) );
  XNOR U11389 ( .A(n11566), .B(n11570), .Z(n11568) );
  XOR U11390 ( .A(n11451), .B(n11571), .Z(n11444) );
  IV U11391 ( .A(n11450), .Z(n11571) );
  XNOR U11392 ( .A(n11447), .B(n11572), .Z(n11450) );
  XOR U11393 ( .A(n11573), .B(n11574), .Z(n11447) );
  ANDN U11394 ( .A(n11575), .B(n11576), .Z(n11574) );
  XNOR U11395 ( .A(n11573), .B(n11577), .Z(n11575) );
  XOR U11396 ( .A(n11458), .B(n11578), .Z(n11451) );
  IV U11397 ( .A(n11457), .Z(n11578) );
  XNOR U11398 ( .A(n11454), .B(n11579), .Z(n11457) );
  XOR U11399 ( .A(n11580), .B(n11581), .Z(n11454) );
  ANDN U11400 ( .A(n11582), .B(n11583), .Z(n11581) );
  XNOR U11401 ( .A(n11580), .B(n11584), .Z(n11582) );
  XOR U11402 ( .A(n11465), .B(n11585), .Z(n11458) );
  IV U11403 ( .A(n11464), .Z(n11585) );
  XNOR U11404 ( .A(n11461), .B(n11586), .Z(n11464) );
  XOR U11405 ( .A(n11587), .B(n11588), .Z(n11461) );
  ANDN U11406 ( .A(n11589), .B(n11590), .Z(n11588) );
  XNOR U11407 ( .A(n11587), .B(n11591), .Z(n11589) );
  XOR U11408 ( .A(n11472), .B(n11592), .Z(n11465) );
  IV U11409 ( .A(n11471), .Z(n11592) );
  XNOR U11410 ( .A(n11468), .B(n11593), .Z(n11471) );
  XOR U11411 ( .A(n11594), .B(n11595), .Z(n11468) );
  ANDN U11412 ( .A(n11596), .B(n11597), .Z(n11595) );
  XNOR U11413 ( .A(n11594), .B(n11598), .Z(n11596) );
  XOR U11414 ( .A(n11479), .B(n11599), .Z(n11472) );
  IV U11415 ( .A(n11478), .Z(n11599) );
  XNOR U11416 ( .A(n11475), .B(n11600), .Z(n11478) );
  XOR U11417 ( .A(n11601), .B(n11602), .Z(n11475) );
  ANDN U11418 ( .A(n11603), .B(n11604), .Z(n11602) );
  XNOR U11419 ( .A(n11601), .B(n11605), .Z(n11603) );
  XOR U11420 ( .A(n11485), .B(n11606), .Z(n11479) );
  IV U11421 ( .A(n11484), .Z(n11606) );
  XNOR U11422 ( .A(n11481), .B(n11607), .Z(n11484) );
  XOR U11423 ( .A(n11608), .B(n11609), .Z(n11481) );
  ANDN U11424 ( .A(n11610), .B(n11611), .Z(n11609) );
  XNOR U11425 ( .A(n11608), .B(n11612), .Z(n11610) );
  XOR U11426 ( .A(n11491), .B(n11613), .Z(n11485) );
  IV U11427 ( .A(n11490), .Z(n11613) );
  XNOR U11428 ( .A(n11487), .B(n11600), .Z(n11490) );
  AND U11429 ( .A(n11869), .B(n11341), .Z(n11600) );
  XOR U11430 ( .A(n11614), .B(n11615), .Z(n11487) );
  ANDN U11431 ( .A(n11616), .B(n11617), .Z(n11615) );
  XNOR U11432 ( .A(n11614), .B(n11618), .Z(n11616) );
  XOR U11433 ( .A(n11497), .B(n11619), .Z(n11491) );
  IV U11434 ( .A(n11496), .Z(n11619) );
  XNOR U11435 ( .A(n11493), .B(n11593), .Z(n11496) );
  AND U11436 ( .A(n12128), .B(n11049), .Z(n11593) );
  XOR U11437 ( .A(n11620), .B(n11621), .Z(n11493) );
  ANDN U11438 ( .A(n11622), .B(n11623), .Z(n11621) );
  XNOR U11439 ( .A(n11620), .B(n11624), .Z(n11622) );
  XOR U11440 ( .A(n11503), .B(n11625), .Z(n11497) );
  IV U11441 ( .A(n11502), .Z(n11625) );
  XNOR U11442 ( .A(n11499), .B(n11586), .Z(n11502) );
  AND U11443 ( .A(n12387), .B(n10731), .Z(n11586) );
  XOR U11444 ( .A(n11626), .B(n11627), .Z(n11499) );
  ANDN U11445 ( .A(n11628), .B(n11629), .Z(n11627) );
  XNOR U11446 ( .A(n11626), .B(n11630), .Z(n11628) );
  XOR U11447 ( .A(n11509), .B(n11631), .Z(n11503) );
  IV U11448 ( .A(n11508), .Z(n11631) );
  XNOR U11449 ( .A(n11505), .B(n11579), .Z(n11508) );
  AND U11450 ( .A(n12644), .B(n10387), .Z(n11579) );
  XOR U11451 ( .A(n11632), .B(n11633), .Z(n11505) );
  ANDN U11452 ( .A(n11634), .B(n11635), .Z(n11633) );
  XNOR U11453 ( .A(n11632), .B(n11636), .Z(n11634) );
  XOR U11454 ( .A(n11515), .B(n11637), .Z(n11509) );
  IV U11455 ( .A(n11514), .Z(n11637) );
  XNOR U11456 ( .A(n11511), .B(n11572), .Z(n11514) );
  AND U11457 ( .A(n12880), .B(n10017), .Z(n11572) );
  XOR U11458 ( .A(n11638), .B(n11639), .Z(n11511) );
  ANDN U11459 ( .A(n11640), .B(n11641), .Z(n11639) );
  XNOR U11460 ( .A(n11638), .B(n11642), .Z(n11640) );
  XOR U11461 ( .A(n11521), .B(n11643), .Z(n11515) );
  IV U11462 ( .A(n11520), .Z(n11643) );
  XNOR U11463 ( .A(n11517), .B(n11565), .Z(n11520) );
  AND U11464 ( .A(n13070), .B(n9621), .Z(n11565) );
  XOR U11465 ( .A(n11644), .B(n11645), .Z(n11517) );
  ANDN U11466 ( .A(n11646), .B(n11647), .Z(n11645) );
  XNOR U11467 ( .A(n11644), .B(n11648), .Z(n11646) );
  XOR U11468 ( .A(n11527), .B(n11649), .Z(n11521) );
  IV U11469 ( .A(n11526), .Z(n11649) );
  XNOR U11470 ( .A(n11523), .B(n11558), .Z(n11526) );
  AND U11471 ( .A(n13207), .B(n9198), .Z(n11558) );
  XOR U11472 ( .A(n11650), .B(n11651), .Z(n11523) );
  ANDN U11473 ( .A(n11652), .B(n11653), .Z(n11651) );
  XNOR U11474 ( .A(n11650), .B(n11654), .Z(n11652) );
  XNOR U11475 ( .A(n11532), .B(n11422), .Z(n11527) );
  XNOR U11476 ( .A(n11529), .B(n11655), .Z(n11532) );
  AND U11477 ( .A(n6527), .B(n8748), .Z(n11655) );
  XOR U11478 ( .A(n11656), .B(n11657), .Z(n11529) );
  ANDN U11479 ( .A(n11658), .B(n11659), .Z(n11657) );
  XNOR U11480 ( .A(n11555), .B(n11656), .Z(n11658) );
  XOR U11481 ( .A(n11660), .B(n11422), .Z(n11552) );
  NANDN U11482 ( .B(n6808), .A(n8272), .Z(n11422) );
  XOR U11483 ( .A(n11661), .B(n11662), .Z(n8272) );
  AND U11484 ( .A(n6809), .B(n11663), .Z(n11662) );
  XNOR U11485 ( .A(n11661), .B(n11539), .Z(n11663) );
  XOR U11486 ( .A(n11537), .B(n11661), .Z(n11539) );
  XOR U11487 ( .A(n11664), .B(n11665), .Z(n11537) );
  ANDN U11488 ( .A(n11664), .B(n11666), .Z(n11665) );
  XOR U11489 ( .A(n11667), .B(n7368), .Z(n11661) );
  IV U11490 ( .A(n11541), .Z(n11660) );
  XOR U11491 ( .A(n11668), .B(n11669), .Z(n11541) );
  AND U11492 ( .A(n11670), .B(n11671), .Z(n11669) );
  XNOR U11493 ( .A(n11668), .B(n11672), .Z(n11671) );
  XNOR U11494 ( .A(n11545), .B(n11548), .Z(n11551) );
  XOR U11495 ( .A(n11673), .B(n11674), .Z(n11545) );
  XOR U11496 ( .A(n11675), .B(n11676), .Z(n11548) );
  AND U11497 ( .A(n11677), .B(n11678), .Z(n11676) );
  XOR U11498 ( .A(n11675), .B(n11679), .Z(n11678) );
  XOR U11499 ( .A(n11680), .B(n11681), .Z(n11679) );
  ANDN U11500 ( .A(n11682), .B(n11683), .Z(n11680) );
  XOR U11501 ( .A(n11684), .B(n11681), .Z(n11682) );
  XOR U11502 ( .A(n11685), .B(n11672), .Z(n11677) );
  XOR U11503 ( .A(n11686), .B(n11687), .Z(n11672) );
  XNOR U11504 ( .A(n11670), .B(n11675), .Z(n11685) );
  XOR U11505 ( .A(n11688), .B(n11556), .Z(n11670) );
  XOR U11506 ( .A(n11563), .B(n11689), .Z(n11556) );
  IV U11507 ( .A(n11561), .Z(n11689) );
  XNOR U11508 ( .A(n11690), .B(n11560), .Z(n11561) );
  OR U11509 ( .A(n11691), .B(n11692), .Z(n11560) );
  NANDN U11510 ( .B(n6541), .A(n9198), .Z(n11690) );
  XOR U11511 ( .A(n11570), .B(n11693), .Z(n11563) );
  IV U11512 ( .A(n11569), .Z(n11693) );
  XNOR U11513 ( .A(n11566), .B(n11694), .Z(n11569) );
  XOR U11514 ( .A(n11695), .B(n11696), .Z(n11566) );
  NANDN U11515 ( .B(n11697), .A(n11698), .Z(n11695) );
  XOR U11516 ( .A(n11696), .B(n11699), .Z(n11698) );
  XOR U11517 ( .A(n11577), .B(n11700), .Z(n11570) );
  IV U11518 ( .A(n11576), .Z(n11700) );
  XNOR U11519 ( .A(n11573), .B(n11701), .Z(n11576) );
  XOR U11520 ( .A(n11702), .B(n11703), .Z(n11573) );
  ANDN U11521 ( .A(n11704), .B(n11705), .Z(n11703) );
  XNOR U11522 ( .A(n11702), .B(n11706), .Z(n11704) );
  XOR U11523 ( .A(n11584), .B(n11707), .Z(n11577) );
  IV U11524 ( .A(n11583), .Z(n11707) );
  XNOR U11525 ( .A(n11580), .B(n11708), .Z(n11583) );
  XOR U11526 ( .A(n11709), .B(n11710), .Z(n11580) );
  ANDN U11527 ( .A(n11711), .B(n11712), .Z(n11710) );
  XNOR U11528 ( .A(n11709), .B(n11713), .Z(n11711) );
  XOR U11529 ( .A(n11591), .B(n11714), .Z(n11584) );
  IV U11530 ( .A(n11590), .Z(n11714) );
  XNOR U11531 ( .A(n11587), .B(n11715), .Z(n11590) );
  XOR U11532 ( .A(n11716), .B(n11717), .Z(n11587) );
  ANDN U11533 ( .A(n11718), .B(n11719), .Z(n11717) );
  XNOR U11534 ( .A(n11716), .B(n11720), .Z(n11718) );
  XOR U11535 ( .A(n11598), .B(n11721), .Z(n11591) );
  IV U11536 ( .A(n11597), .Z(n11721) );
  XNOR U11537 ( .A(n11594), .B(n11722), .Z(n11597) );
  XOR U11538 ( .A(n11723), .B(n11724), .Z(n11594) );
  ANDN U11539 ( .A(n11725), .B(n11726), .Z(n11724) );
  XNOR U11540 ( .A(n11723), .B(n11727), .Z(n11725) );
  XOR U11541 ( .A(n11605), .B(n11728), .Z(n11598) );
  IV U11542 ( .A(n11604), .Z(n11728) );
  XNOR U11543 ( .A(n11601), .B(n11729), .Z(n11604) );
  XOR U11544 ( .A(n11730), .B(n11731), .Z(n11601) );
  ANDN U11545 ( .A(n11732), .B(n11733), .Z(n11731) );
  XNOR U11546 ( .A(n11730), .B(n11734), .Z(n11732) );
  XOR U11547 ( .A(n11612), .B(n11735), .Z(n11605) );
  IV U11548 ( .A(n11611), .Z(n11735) );
  XNOR U11549 ( .A(n11608), .B(n11736), .Z(n11611) );
  XOR U11550 ( .A(n11737), .B(n11738), .Z(n11608) );
  ANDN U11551 ( .A(n11739), .B(n11740), .Z(n11738) );
  XNOR U11552 ( .A(n11737), .B(n11741), .Z(n11739) );
  XOR U11553 ( .A(n11618), .B(n11742), .Z(n11612) );
  IV U11554 ( .A(n11617), .Z(n11742) );
  XNOR U11555 ( .A(n11614), .B(n11736), .Z(n11617) );
  AND U11556 ( .A(n11869), .B(n11607), .Z(n11736) );
  XOR U11557 ( .A(n11743), .B(n11744), .Z(n11614) );
  ANDN U11558 ( .A(n11745), .B(n11746), .Z(n11744) );
  XNOR U11559 ( .A(n11743), .B(n11747), .Z(n11745) );
  XOR U11560 ( .A(n11624), .B(n11748), .Z(n11618) );
  IV U11561 ( .A(n11623), .Z(n11748) );
  XNOR U11562 ( .A(n11620), .B(n11729), .Z(n11623) );
  AND U11563 ( .A(n12128), .B(n11341), .Z(n11729) );
  XOR U11564 ( .A(n11749), .B(n11750), .Z(n11620) );
  ANDN U11565 ( .A(n11751), .B(n11752), .Z(n11750) );
  XNOR U11566 ( .A(n11749), .B(n11753), .Z(n11751) );
  XOR U11567 ( .A(n11630), .B(n11754), .Z(n11624) );
  IV U11568 ( .A(n11629), .Z(n11754) );
  XNOR U11569 ( .A(n11626), .B(n11722), .Z(n11629) );
  AND U11570 ( .A(n12387), .B(n11049), .Z(n11722) );
  XOR U11571 ( .A(n11755), .B(n11756), .Z(n11626) );
  ANDN U11572 ( .A(n11757), .B(n11758), .Z(n11756) );
  XNOR U11573 ( .A(n11755), .B(n11759), .Z(n11757) );
  XOR U11574 ( .A(n11636), .B(n11760), .Z(n11630) );
  IV U11575 ( .A(n11635), .Z(n11760) );
  XNOR U11576 ( .A(n11632), .B(n11715), .Z(n11635) );
  AND U11577 ( .A(n12644), .B(n10731), .Z(n11715) );
  XOR U11578 ( .A(n11761), .B(n11762), .Z(n11632) );
  ANDN U11579 ( .A(n11763), .B(n11764), .Z(n11762) );
  XNOR U11580 ( .A(n11761), .B(n11765), .Z(n11763) );
  XOR U11581 ( .A(n11642), .B(n11766), .Z(n11636) );
  IV U11582 ( .A(n11641), .Z(n11766) );
  XNOR U11583 ( .A(n11638), .B(n11708), .Z(n11641) );
  AND U11584 ( .A(n12880), .B(n10387), .Z(n11708) );
  XOR U11585 ( .A(n11767), .B(n11768), .Z(n11638) );
  ANDN U11586 ( .A(n11769), .B(n11770), .Z(n11768) );
  XNOR U11587 ( .A(n11767), .B(n11771), .Z(n11769) );
  XOR U11588 ( .A(n11648), .B(n11772), .Z(n11642) );
  IV U11589 ( .A(n11647), .Z(n11772) );
  XNOR U11590 ( .A(n11644), .B(n11701), .Z(n11647) );
  AND U11591 ( .A(n13070), .B(n10017), .Z(n11701) );
  XOR U11592 ( .A(n11773), .B(n11774), .Z(n11644) );
  ANDN U11593 ( .A(n11775), .B(n11776), .Z(n11774) );
  XNOR U11594 ( .A(n11773), .B(n11777), .Z(n11775) );
  XOR U11595 ( .A(n11654), .B(n11778), .Z(n11648) );
  IV U11596 ( .A(n11653), .Z(n11778) );
  XNOR U11597 ( .A(n11650), .B(n11694), .Z(n11653) );
  AND U11598 ( .A(n13207), .B(n9621), .Z(n11694) );
  XOR U11599 ( .A(n11779), .B(n11780), .Z(n11650) );
  ANDN U11600 ( .A(n11781), .B(n11782), .Z(n11780) );
  XNOR U11601 ( .A(n11779), .B(n11783), .Z(n11781) );
  XNOR U11602 ( .A(n11659), .B(n11555), .Z(n11654) );
  XNOR U11603 ( .A(n11656), .B(n11784), .Z(n11659) );
  AND U11604 ( .A(n6527), .B(n9198), .Z(n11784) );
  XOR U11605 ( .A(n11785), .B(n11786), .Z(n11656) );
  ANDN U11606 ( .A(n11787), .B(n11788), .Z(n11786) );
  XNOR U11607 ( .A(n11691), .B(n11785), .Z(n11787) );
  XOR U11608 ( .A(n11789), .B(n11555), .Z(n11688) );
  NANDN U11609 ( .B(n6808), .A(n8748), .Z(n11555) );
  XOR U11610 ( .A(n11790), .B(n11791), .Z(n8748) );
  AND U11611 ( .A(n6809), .B(n11792), .Z(n11791) );
  XNOR U11612 ( .A(n11790), .B(n11666), .Z(n11792) );
  XOR U11613 ( .A(n11664), .B(n11790), .Z(n11666) );
  XOR U11614 ( .A(n11793), .B(n11794), .Z(n11664) );
  ANDN U11615 ( .A(n11793), .B(n11795), .Z(n11794) );
  XOR U11616 ( .A(n11796), .B(n7368), .Z(n11790) );
  IV U11617 ( .A(n11668), .Z(n11789) );
  XOR U11618 ( .A(n11797), .B(n11798), .Z(n11668) );
  AND U11619 ( .A(n11799), .B(n11800), .Z(n11798) );
  XNOR U11620 ( .A(n11797), .B(n11801), .Z(n11800) );
  XOR U11621 ( .A(n11802), .B(n11803), .Z(n11675) );
  AND U11622 ( .A(n11804), .B(n11805), .Z(n11803) );
  XNOR U11623 ( .A(n11683), .B(n11806), .Z(n11805) );
  XOR U11624 ( .A(n11802), .B(n11684), .Z(n11806) );
  XOR U11625 ( .A(n11807), .B(n11808), .Z(n11684) );
  ANDN U11626 ( .A(n11809), .B(n11810), .Z(n11808) );
  XNOR U11627 ( .A(n11807), .B(n11811), .Z(n11809) );
  XNOR U11628 ( .A(n11681), .B(n11812), .Z(n11683) );
  XOR U11629 ( .A(n11813), .B(n11814), .Z(n11681) );
  AND U11630 ( .A(n11815), .B(n11816), .Z(n11814) );
  XNOR U11631 ( .A(n11817), .B(n11813), .Z(n11816) );
  XOR U11632 ( .A(n11818), .B(n11801), .Z(n11804) );
  XOR U11633 ( .A(n11819), .B(n11820), .Z(n11801) );
  XNOR U11634 ( .A(n11799), .B(n11802), .Z(n11818) );
  XOR U11635 ( .A(n11821), .B(n11692), .Z(n11799) );
  XOR U11636 ( .A(n11699), .B(n11822), .Z(n11692) );
  IV U11637 ( .A(n11697), .Z(n11822) );
  XNOR U11638 ( .A(n11823), .B(n11696), .Z(n11697) );
  OR U11639 ( .A(n11824), .B(n11825), .Z(n11696) );
  NANDN U11640 ( .B(n6541), .A(n9621), .Z(n11823) );
  XOR U11641 ( .A(n11706), .B(n11826), .Z(n11699) );
  IV U11642 ( .A(n11705), .Z(n11826) );
  XNOR U11643 ( .A(n11702), .B(n11827), .Z(n11705) );
  XOR U11644 ( .A(n11828), .B(n11829), .Z(n11702) );
  NANDN U11645 ( .B(n11830), .A(n11831), .Z(n11828) );
  XOR U11646 ( .A(n11829), .B(n11832), .Z(n11831) );
  XOR U11647 ( .A(n11713), .B(n11833), .Z(n11706) );
  IV U11648 ( .A(n11712), .Z(n11833) );
  XNOR U11649 ( .A(n11709), .B(n11834), .Z(n11712) );
  XOR U11650 ( .A(n11835), .B(n11836), .Z(n11709) );
  ANDN U11651 ( .A(n11837), .B(n11838), .Z(n11836) );
  XNOR U11652 ( .A(n11835), .B(n11839), .Z(n11837) );
  XOR U11653 ( .A(n11720), .B(n11840), .Z(n11713) );
  IV U11654 ( .A(n11719), .Z(n11840) );
  XNOR U11655 ( .A(n11716), .B(n11841), .Z(n11719) );
  XOR U11656 ( .A(n11842), .B(n11843), .Z(n11716) );
  ANDN U11657 ( .A(n11844), .B(n11845), .Z(n11843) );
  XNOR U11658 ( .A(n11842), .B(n11846), .Z(n11844) );
  XOR U11659 ( .A(n11727), .B(n11847), .Z(n11720) );
  IV U11660 ( .A(n11726), .Z(n11847) );
  XNOR U11661 ( .A(n11723), .B(n11848), .Z(n11726) );
  XOR U11662 ( .A(n11849), .B(n11850), .Z(n11723) );
  ANDN U11663 ( .A(n11851), .B(n11852), .Z(n11850) );
  XNOR U11664 ( .A(n11849), .B(n11853), .Z(n11851) );
  XOR U11665 ( .A(n11734), .B(n11854), .Z(n11727) );
  IV U11666 ( .A(n11733), .Z(n11854) );
  XNOR U11667 ( .A(n11730), .B(n11855), .Z(n11733) );
  XOR U11668 ( .A(n11856), .B(n11857), .Z(n11730) );
  ANDN U11669 ( .A(n11858), .B(n11859), .Z(n11857) );
  XNOR U11670 ( .A(n11856), .B(n11860), .Z(n11858) );
  XOR U11671 ( .A(n11741), .B(n11861), .Z(n11734) );
  IV U11672 ( .A(n11740), .Z(n11861) );
  XNOR U11673 ( .A(n11737), .B(n11862), .Z(n11740) );
  XOR U11674 ( .A(n11863), .B(n11864), .Z(n11737) );
  ANDN U11675 ( .A(n11865), .B(n11866), .Z(n11864) );
  XNOR U11676 ( .A(n11863), .B(n11867), .Z(n11865) );
  XOR U11677 ( .A(n11747), .B(n11868), .Z(n11741) );
  IV U11678 ( .A(n11746), .Z(n11868) );
  XNOR U11679 ( .A(n11743), .B(n11869), .Z(n11746) );
  XOR U11680 ( .A(n11870), .B(n11871), .Z(n11743) );
  ANDN U11681 ( .A(n11872), .B(n11873), .Z(n11871) );
  XNOR U11682 ( .A(n11870), .B(n11874), .Z(n11872) );
  XOR U11683 ( .A(n11753), .B(n11875), .Z(n11747) );
  IV U11684 ( .A(n11752), .Z(n11875) );
  XNOR U11685 ( .A(n11749), .B(n11862), .Z(n11752) );
  AND U11686 ( .A(n12128), .B(n11607), .Z(n11862) );
  XOR U11687 ( .A(n11876), .B(n11877), .Z(n11749) );
  ANDN U11688 ( .A(n11878), .B(n11879), .Z(n11877) );
  XNOR U11689 ( .A(n11876), .B(n11880), .Z(n11878) );
  XOR U11690 ( .A(n11759), .B(n11881), .Z(n11753) );
  IV U11691 ( .A(n11758), .Z(n11881) );
  XNOR U11692 ( .A(n11755), .B(n11855), .Z(n11758) );
  AND U11693 ( .A(n12387), .B(n11341), .Z(n11855) );
  XOR U11694 ( .A(n11882), .B(n11883), .Z(n11755) );
  ANDN U11695 ( .A(n11884), .B(n11885), .Z(n11883) );
  XNOR U11696 ( .A(n11882), .B(n11886), .Z(n11884) );
  XOR U11697 ( .A(n11765), .B(n11887), .Z(n11759) );
  IV U11698 ( .A(n11764), .Z(n11887) );
  XNOR U11699 ( .A(n11761), .B(n11848), .Z(n11764) );
  AND U11700 ( .A(n12644), .B(n11049), .Z(n11848) );
  XOR U11701 ( .A(n11888), .B(n11889), .Z(n11761) );
  ANDN U11702 ( .A(n11890), .B(n11891), .Z(n11889) );
  XNOR U11703 ( .A(n11888), .B(n11892), .Z(n11890) );
  XOR U11704 ( .A(n11771), .B(n11893), .Z(n11765) );
  IV U11705 ( .A(n11770), .Z(n11893) );
  XNOR U11706 ( .A(n11767), .B(n11841), .Z(n11770) );
  AND U11707 ( .A(n12880), .B(n10731), .Z(n11841) );
  XOR U11708 ( .A(n11894), .B(n11895), .Z(n11767) );
  ANDN U11709 ( .A(n11896), .B(n11897), .Z(n11895) );
  XNOR U11710 ( .A(n11894), .B(n11898), .Z(n11896) );
  XOR U11711 ( .A(n11777), .B(n11899), .Z(n11771) );
  IV U11712 ( .A(n11776), .Z(n11899) );
  XNOR U11713 ( .A(n11773), .B(n11834), .Z(n11776) );
  AND U11714 ( .A(n13070), .B(n10387), .Z(n11834) );
  XOR U11715 ( .A(n11900), .B(n11901), .Z(n11773) );
  ANDN U11716 ( .A(n11902), .B(n11903), .Z(n11901) );
  XNOR U11717 ( .A(n11900), .B(n11904), .Z(n11902) );
  XOR U11718 ( .A(n11783), .B(n11905), .Z(n11777) );
  IV U11719 ( .A(n11782), .Z(n11905) );
  XNOR U11720 ( .A(n11779), .B(n11827), .Z(n11782) );
  AND U11721 ( .A(n13207), .B(n10017), .Z(n11827) );
  XOR U11722 ( .A(n11906), .B(n11907), .Z(n11779) );
  ANDN U11723 ( .A(n11908), .B(n11909), .Z(n11907) );
  XNOR U11724 ( .A(n11906), .B(n11910), .Z(n11908) );
  XNOR U11725 ( .A(n11788), .B(n11691), .Z(n11783) );
  XNOR U11726 ( .A(n11785), .B(n11911), .Z(n11788) );
  AND U11727 ( .A(n6527), .B(n9621), .Z(n11911) );
  XOR U11728 ( .A(n11912), .B(n11913), .Z(n11785) );
  ANDN U11729 ( .A(n11914), .B(n11915), .Z(n11913) );
  XNOR U11730 ( .A(n11824), .B(n11912), .Z(n11914) );
  XOR U11731 ( .A(n11916), .B(n11691), .Z(n11821) );
  NANDN U11732 ( .B(n6808), .A(n9198), .Z(n11691) );
  XOR U11733 ( .A(n11917), .B(n11918), .Z(n9198) );
  AND U11734 ( .A(n6809), .B(n11919), .Z(n11918) );
  XNOR U11735 ( .A(n11917), .B(n11795), .Z(n11919) );
  XOR U11736 ( .A(n11793), .B(n11917), .Z(n11795) );
  XOR U11737 ( .A(n11920), .B(n11921), .Z(n11793) );
  ANDN U11738 ( .A(n11920), .B(n11922), .Z(n11921) );
  XOR U11739 ( .A(n11923), .B(n7368), .Z(n11917) );
  IV U11740 ( .A(n11797), .Z(n11916) );
  XOR U11741 ( .A(n11924), .B(n11925), .Z(n11797) );
  AND U11742 ( .A(n11926), .B(n11927), .Z(n11925) );
  XNOR U11743 ( .A(n11924), .B(n11928), .Z(n11927) );
  XOR U11744 ( .A(n11929), .B(n11930), .Z(n11802) );
  AND U11745 ( .A(n11931), .B(n11932), .Z(n11930) );
  XOR U11746 ( .A(n11815), .B(n11933), .Z(n11932) );
  XNOR U11747 ( .A(n11929), .B(n11817), .Z(n11933) );
  XOR U11748 ( .A(n11811), .B(n11934), .Z(n11817) );
  IV U11749 ( .A(n11810), .Z(n11934) );
  XNOR U11750 ( .A(n11807), .B(n11935), .Z(n11810) );
  XOR U11751 ( .A(n11936), .B(n11937), .Z(n11807) );
  ANDN U11752 ( .A(n11938), .B(n11939), .Z(n11937) );
  XNOR U11753 ( .A(n11936), .B(n11940), .Z(n11938) );
  XNOR U11754 ( .A(n11941), .B(n11942), .Z(n11811) );
  ANDN U11755 ( .A(n11943), .B(n11944), .Z(n11942) );
  XNOR U11756 ( .A(n11941), .B(n11945), .Z(n11943) );
  XOR U11757 ( .A(n11813), .B(n11935), .Z(n11815) );
  AND U11758 ( .A(n11812), .B(n12061), .Z(n11935) );
  XOR U11759 ( .A(n11946), .B(n11947), .Z(n11813) );
  AND U11760 ( .A(n11948), .B(n11949), .Z(n11947) );
  XNOR U11761 ( .A(n11950), .B(n11946), .Z(n11949) );
  XOR U11762 ( .A(n11951), .B(n11928), .Z(n11931) );
  XOR U11763 ( .A(n11952), .B(n11953), .Z(n11928) );
  XNOR U11764 ( .A(n11926), .B(n11929), .Z(n11951) );
  XOR U11765 ( .A(n11954), .B(n11825), .Z(n11926) );
  XOR U11766 ( .A(n11832), .B(n11955), .Z(n11825) );
  IV U11767 ( .A(n11830), .Z(n11955) );
  XNOR U11768 ( .A(n11956), .B(n11829), .Z(n11830) );
  OR U11769 ( .A(n11957), .B(n11958), .Z(n11829) );
  NANDN U11770 ( .B(n6541), .A(n10017), .Z(n11956) );
  XOR U11771 ( .A(n11839), .B(n11959), .Z(n11832) );
  IV U11772 ( .A(n11838), .Z(n11959) );
  XNOR U11773 ( .A(n11835), .B(n11960), .Z(n11838) );
  XOR U11774 ( .A(n11961), .B(n11962), .Z(n11835) );
  NANDN U11775 ( .B(n11963), .A(n11964), .Z(n11961) );
  XOR U11776 ( .A(n11962), .B(n11965), .Z(n11964) );
  XOR U11777 ( .A(n11846), .B(n11966), .Z(n11839) );
  IV U11778 ( .A(n11845), .Z(n11966) );
  XNOR U11779 ( .A(n11842), .B(n11967), .Z(n11845) );
  XOR U11780 ( .A(n11968), .B(n11969), .Z(n11842) );
  ANDN U11781 ( .A(n11970), .B(n11971), .Z(n11969) );
  XNOR U11782 ( .A(n11968), .B(n11972), .Z(n11970) );
  XOR U11783 ( .A(n11853), .B(n11973), .Z(n11846) );
  IV U11784 ( .A(n11852), .Z(n11973) );
  XNOR U11785 ( .A(n11849), .B(n11974), .Z(n11852) );
  XOR U11786 ( .A(n11975), .B(n11976), .Z(n11849) );
  ANDN U11787 ( .A(n11977), .B(n11978), .Z(n11976) );
  XNOR U11788 ( .A(n11975), .B(n11979), .Z(n11977) );
  XOR U11789 ( .A(n11860), .B(n11980), .Z(n11853) );
  IV U11790 ( .A(n11859), .Z(n11980) );
  XNOR U11791 ( .A(n11856), .B(n11981), .Z(n11859) );
  XOR U11792 ( .A(n11982), .B(n11983), .Z(n11856) );
  ANDN U11793 ( .A(n11984), .B(n11985), .Z(n11983) );
  XNOR U11794 ( .A(n11982), .B(n11986), .Z(n11984) );
  XOR U11795 ( .A(n11867), .B(n11987), .Z(n11860) );
  IV U11796 ( .A(n11866), .Z(n11987) );
  XNOR U11797 ( .A(n11863), .B(n11988), .Z(n11866) );
  XOR U11798 ( .A(n11989), .B(n11990), .Z(n11863) );
  ANDN U11799 ( .A(n11991), .B(n11992), .Z(n11990) );
  XNOR U11800 ( .A(n11989), .B(n11993), .Z(n11991) );
  XOR U11801 ( .A(n11874), .B(n11994), .Z(n11867) );
  IV U11802 ( .A(n11873), .Z(n11994) );
  XNOR U11803 ( .A(n11870), .B(n11995), .Z(n11873) );
  XOR U11804 ( .A(n11996), .B(n11997), .Z(n11870) );
  ANDN U11805 ( .A(n11998), .B(n11999), .Z(n11997) );
  XNOR U11806 ( .A(n11996), .B(n12000), .Z(n11998) );
  XOR U11807 ( .A(n11880), .B(n12001), .Z(n11874) );
  IV U11808 ( .A(n11879), .Z(n12001) );
  XNOR U11809 ( .A(n11876), .B(n11995), .Z(n11879) );
  AND U11810 ( .A(n12128), .B(n11869), .Z(n11995) );
  XOR U11811 ( .A(n12002), .B(n12003), .Z(n11876) );
  ANDN U11812 ( .A(n12004), .B(n12005), .Z(n12003) );
  XNOR U11813 ( .A(n12002), .B(n12006), .Z(n12004) );
  XOR U11814 ( .A(n11886), .B(n12007), .Z(n11880) );
  IV U11815 ( .A(n11885), .Z(n12007) );
  XNOR U11816 ( .A(n11882), .B(n11988), .Z(n11885) );
  AND U11817 ( .A(n12387), .B(n11607), .Z(n11988) );
  XOR U11818 ( .A(n12008), .B(n12009), .Z(n11882) );
  ANDN U11819 ( .A(n12010), .B(n12011), .Z(n12009) );
  XNOR U11820 ( .A(n12008), .B(n12012), .Z(n12010) );
  XOR U11821 ( .A(n11892), .B(n12013), .Z(n11886) );
  IV U11822 ( .A(n11891), .Z(n12013) );
  XNOR U11823 ( .A(n11888), .B(n11981), .Z(n11891) );
  AND U11824 ( .A(n12644), .B(n11341), .Z(n11981) );
  XOR U11825 ( .A(n12014), .B(n12015), .Z(n11888) );
  ANDN U11826 ( .A(n12016), .B(n12017), .Z(n12015) );
  XNOR U11827 ( .A(n12014), .B(n12018), .Z(n12016) );
  XOR U11828 ( .A(n11898), .B(n12019), .Z(n11892) );
  IV U11829 ( .A(n11897), .Z(n12019) );
  XNOR U11830 ( .A(n11894), .B(n11974), .Z(n11897) );
  AND U11831 ( .A(n12880), .B(n11049), .Z(n11974) );
  XOR U11832 ( .A(n12020), .B(n12021), .Z(n11894) );
  ANDN U11833 ( .A(n12022), .B(n12023), .Z(n12021) );
  XNOR U11834 ( .A(n12020), .B(n12024), .Z(n12022) );
  XOR U11835 ( .A(n11904), .B(n12025), .Z(n11898) );
  IV U11836 ( .A(n11903), .Z(n12025) );
  XNOR U11837 ( .A(n11900), .B(n11967), .Z(n11903) );
  AND U11838 ( .A(n13070), .B(n10731), .Z(n11967) );
  XOR U11839 ( .A(n12026), .B(n12027), .Z(n11900) );
  ANDN U11840 ( .A(n12028), .B(n12029), .Z(n12027) );
  XNOR U11841 ( .A(n12026), .B(n12030), .Z(n12028) );
  XOR U11842 ( .A(n11910), .B(n12031), .Z(n11904) );
  IV U11843 ( .A(n11909), .Z(n12031) );
  XNOR U11844 ( .A(n11906), .B(n11960), .Z(n11909) );
  AND U11845 ( .A(n13207), .B(n10387), .Z(n11960) );
  XOR U11846 ( .A(n12032), .B(n12033), .Z(n11906) );
  ANDN U11847 ( .A(n12034), .B(n12035), .Z(n12033) );
  XNOR U11848 ( .A(n12032), .B(n12036), .Z(n12034) );
  XNOR U11849 ( .A(n11915), .B(n11824), .Z(n11910) );
  XNOR U11850 ( .A(n11912), .B(n12037), .Z(n11915) );
  AND U11851 ( .A(n6527), .B(n10017), .Z(n12037) );
  XOR U11852 ( .A(n12038), .B(n12039), .Z(n11912) );
  ANDN U11853 ( .A(n12040), .B(n12041), .Z(n12039) );
  XNOR U11854 ( .A(n11957), .B(n12038), .Z(n12040) );
  XOR U11855 ( .A(n12042), .B(n11824), .Z(n11954) );
  NANDN U11856 ( .B(n6808), .A(n9621), .Z(n11824) );
  XOR U11857 ( .A(n12043), .B(n12044), .Z(n9621) );
  AND U11858 ( .A(n6809), .B(n12045), .Z(n12044) );
  XNOR U11859 ( .A(n12043), .B(n11922), .Z(n12045) );
  XOR U11860 ( .A(n11920), .B(n12043), .Z(n11922) );
  XOR U11861 ( .A(n12046), .B(n12047), .Z(n11920) );
  ANDN U11862 ( .A(n12046), .B(n12048), .Z(n12047) );
  XOR U11863 ( .A(n12049), .B(n7368), .Z(n12043) );
  IV U11864 ( .A(n11924), .Z(n12042) );
  XOR U11865 ( .A(n12050), .B(n12051), .Z(n11924) );
  AND U11866 ( .A(n12052), .B(n12053), .Z(n12051) );
  XNOR U11867 ( .A(n12050), .B(n12054), .Z(n12053) );
  XOR U11868 ( .A(n12055), .B(n12056), .Z(n11929) );
  AND U11869 ( .A(n12057), .B(n12058), .Z(n12056) );
  XOR U11870 ( .A(n11948), .B(n12059), .Z(n12058) );
  XNOR U11871 ( .A(n12055), .B(n11950), .Z(n12059) );
  XOR U11872 ( .A(n11940), .B(n12060), .Z(n11950) );
  IV U11873 ( .A(n11939), .Z(n12060) );
  XNOR U11874 ( .A(n11936), .B(n12061), .Z(n11939) );
  XOR U11875 ( .A(n12062), .B(n12063), .Z(n11936) );
  ANDN U11876 ( .A(n12064), .B(n12065), .Z(n12063) );
  XNOR U11877 ( .A(n12062), .B(n12066), .Z(n12064) );
  XOR U11878 ( .A(n11945), .B(n12067), .Z(n11940) );
  IV U11879 ( .A(n11944), .Z(n12067) );
  XNOR U11880 ( .A(n11941), .B(n12068), .Z(n11944) );
  XOR U11881 ( .A(n12069), .B(n12070), .Z(n11941) );
  ANDN U11882 ( .A(n12071), .B(n12072), .Z(n12070) );
  XNOR U11883 ( .A(n12069), .B(n12073), .Z(n12071) );
  XNOR U11884 ( .A(n12074), .B(n12075), .Z(n11945) );
  ANDN U11885 ( .A(n12076), .B(n12077), .Z(n12075) );
  XNOR U11886 ( .A(n12074), .B(n12078), .Z(n12076) );
  XOR U11887 ( .A(n11946), .B(n12068), .Z(n11948) );
  AND U11888 ( .A(n11812), .B(n12321), .Z(n12068) );
  XOR U11889 ( .A(n12079), .B(n12080), .Z(n11946) );
  AND U11890 ( .A(n12081), .B(n12082), .Z(n12080) );
  XNOR U11891 ( .A(n12083), .B(n12079), .Z(n12082) );
  XOR U11892 ( .A(n12084), .B(n12054), .Z(n12057) );
  XOR U11893 ( .A(n12085), .B(n12086), .Z(n12054) );
  XNOR U11894 ( .A(n12052), .B(n12055), .Z(n12084) );
  XOR U11895 ( .A(n12087), .B(n11958), .Z(n12052) );
  XOR U11896 ( .A(n11965), .B(n12088), .Z(n11958) );
  IV U11897 ( .A(n11963), .Z(n12088) );
  XNOR U11898 ( .A(n12089), .B(n11962), .Z(n11963) );
  OR U11899 ( .A(n12090), .B(n12091), .Z(n11962) );
  NANDN U11900 ( .B(n6541), .A(n10387), .Z(n12089) );
  XOR U11901 ( .A(n11972), .B(n12092), .Z(n11965) );
  IV U11902 ( .A(n11971), .Z(n12092) );
  XNOR U11903 ( .A(n11968), .B(n12093), .Z(n11971) );
  XOR U11904 ( .A(n12094), .B(n12095), .Z(n11968) );
  NANDN U11905 ( .B(n12096), .A(n12097), .Z(n12094) );
  XOR U11906 ( .A(n12095), .B(n12098), .Z(n12097) );
  XOR U11907 ( .A(n11979), .B(n12099), .Z(n11972) );
  IV U11908 ( .A(n11978), .Z(n12099) );
  XNOR U11909 ( .A(n11975), .B(n12100), .Z(n11978) );
  XOR U11910 ( .A(n12101), .B(n12102), .Z(n11975) );
  ANDN U11911 ( .A(n12103), .B(n12104), .Z(n12102) );
  XNOR U11912 ( .A(n12101), .B(n12105), .Z(n12103) );
  XOR U11913 ( .A(n11986), .B(n12106), .Z(n11979) );
  IV U11914 ( .A(n11985), .Z(n12106) );
  XNOR U11915 ( .A(n11982), .B(n12107), .Z(n11985) );
  XOR U11916 ( .A(n12108), .B(n12109), .Z(n11982) );
  ANDN U11917 ( .A(n12110), .B(n12111), .Z(n12109) );
  XNOR U11918 ( .A(n12108), .B(n12112), .Z(n12110) );
  XOR U11919 ( .A(n11993), .B(n12113), .Z(n11986) );
  IV U11920 ( .A(n11992), .Z(n12113) );
  XNOR U11921 ( .A(n11989), .B(n12114), .Z(n11992) );
  XOR U11922 ( .A(n12115), .B(n12116), .Z(n11989) );
  ANDN U11923 ( .A(n12117), .B(n12118), .Z(n12116) );
  XNOR U11924 ( .A(n12115), .B(n12119), .Z(n12117) );
  XOR U11925 ( .A(n12000), .B(n12120), .Z(n11993) );
  IV U11926 ( .A(n11999), .Z(n12120) );
  XNOR U11927 ( .A(n11996), .B(n12121), .Z(n11999) );
  XOR U11928 ( .A(n12122), .B(n12123), .Z(n11996) );
  ANDN U11929 ( .A(n12124), .B(n12125), .Z(n12123) );
  XNOR U11930 ( .A(n12122), .B(n12126), .Z(n12124) );
  XOR U11931 ( .A(n12006), .B(n12127), .Z(n12000) );
  IV U11932 ( .A(n12005), .Z(n12127) );
  XNOR U11933 ( .A(n12002), .B(n12128), .Z(n12005) );
  XOR U11934 ( .A(n12129), .B(n12130), .Z(n12002) );
  ANDN U11935 ( .A(n12131), .B(n12132), .Z(n12130) );
  XNOR U11936 ( .A(n12129), .B(n12133), .Z(n12131) );
  XOR U11937 ( .A(n12012), .B(n12134), .Z(n12006) );
  IV U11938 ( .A(n12011), .Z(n12134) );
  XNOR U11939 ( .A(n12008), .B(n12121), .Z(n12011) );
  AND U11940 ( .A(n12387), .B(n11869), .Z(n12121) );
  XOR U11941 ( .A(n12135), .B(n12136), .Z(n12008) );
  ANDN U11942 ( .A(n12137), .B(n12138), .Z(n12136) );
  XNOR U11943 ( .A(n12135), .B(n12139), .Z(n12137) );
  XOR U11944 ( .A(n12018), .B(n12140), .Z(n12012) );
  IV U11945 ( .A(n12017), .Z(n12140) );
  XNOR U11946 ( .A(n12014), .B(n12114), .Z(n12017) );
  AND U11947 ( .A(n12644), .B(n11607), .Z(n12114) );
  XOR U11948 ( .A(n12141), .B(n12142), .Z(n12014) );
  ANDN U11949 ( .A(n12143), .B(n12144), .Z(n12142) );
  XNOR U11950 ( .A(n12141), .B(n12145), .Z(n12143) );
  XOR U11951 ( .A(n12024), .B(n12146), .Z(n12018) );
  IV U11952 ( .A(n12023), .Z(n12146) );
  XNOR U11953 ( .A(n12020), .B(n12107), .Z(n12023) );
  AND U11954 ( .A(n12880), .B(n11341), .Z(n12107) );
  XOR U11955 ( .A(n12147), .B(n12148), .Z(n12020) );
  ANDN U11956 ( .A(n12149), .B(n12150), .Z(n12148) );
  XNOR U11957 ( .A(n12147), .B(n12151), .Z(n12149) );
  XOR U11958 ( .A(n12030), .B(n12152), .Z(n12024) );
  IV U11959 ( .A(n12029), .Z(n12152) );
  XNOR U11960 ( .A(n12026), .B(n12100), .Z(n12029) );
  AND U11961 ( .A(n13070), .B(n11049), .Z(n12100) );
  XOR U11962 ( .A(n12153), .B(n12154), .Z(n12026) );
  ANDN U11963 ( .A(n12155), .B(n12156), .Z(n12154) );
  XNOR U11964 ( .A(n12153), .B(n12157), .Z(n12155) );
  XOR U11965 ( .A(n12036), .B(n12158), .Z(n12030) );
  IV U11966 ( .A(n12035), .Z(n12158) );
  XNOR U11967 ( .A(n12032), .B(n12093), .Z(n12035) );
  AND U11968 ( .A(n13207), .B(n10731), .Z(n12093) );
  XOR U11969 ( .A(n12159), .B(n12160), .Z(n12032) );
  ANDN U11970 ( .A(n12161), .B(n12162), .Z(n12160) );
  XNOR U11971 ( .A(n12159), .B(n12163), .Z(n12161) );
  XNOR U11972 ( .A(n12041), .B(n11957), .Z(n12036) );
  XNOR U11973 ( .A(n12038), .B(n12164), .Z(n12041) );
  AND U11974 ( .A(n6527), .B(n10387), .Z(n12164) );
  XOR U11975 ( .A(n12165), .B(n12166), .Z(n12038) );
  ANDN U11976 ( .A(n12167), .B(n12168), .Z(n12166) );
  XNOR U11977 ( .A(n12090), .B(n12165), .Z(n12167) );
  XOR U11978 ( .A(n12169), .B(n11957), .Z(n12087) );
  NANDN U11979 ( .B(n6808), .A(n10017), .Z(n11957) );
  XOR U11980 ( .A(n12170), .B(n12171), .Z(n10017) );
  AND U11981 ( .A(n6809), .B(n12172), .Z(n12171) );
  XNOR U11982 ( .A(n12170), .B(n12048), .Z(n12172) );
  XOR U11983 ( .A(n12046), .B(n12170), .Z(n12048) );
  XOR U11984 ( .A(n12173), .B(n12174), .Z(n12046) );
  ANDN U11985 ( .A(n12173), .B(n12175), .Z(n12174) );
  XOR U11986 ( .A(n12176), .B(n7368), .Z(n12170) );
  IV U11987 ( .A(n12050), .Z(n12169) );
  XOR U11988 ( .A(n12177), .B(n12178), .Z(n12050) );
  AND U11989 ( .A(n12179), .B(n12180), .Z(n12178) );
  XNOR U11990 ( .A(n12177), .B(n12181), .Z(n12180) );
  XOR U11991 ( .A(n12182), .B(n12183), .Z(n12055) );
  AND U11992 ( .A(n12184), .B(n12185), .Z(n12183) );
  XOR U11993 ( .A(n12081), .B(n12186), .Z(n12185) );
  XNOR U11994 ( .A(n12182), .B(n12083), .Z(n12186) );
  XOR U11995 ( .A(n12066), .B(n12187), .Z(n12083) );
  IV U11996 ( .A(n12065), .Z(n12187) );
  XNOR U11997 ( .A(n12062), .B(n12188), .Z(n12065) );
  XOR U11998 ( .A(n12189), .B(n12190), .Z(n12062) );
  ANDN U11999 ( .A(n12191), .B(n12192), .Z(n12190) );
  XNOR U12000 ( .A(n12189), .B(n12193), .Z(n12191) );
  XOR U12001 ( .A(n12073), .B(n12194), .Z(n12066) );
  IV U12002 ( .A(n12072), .Z(n12194) );
  XNOR U12003 ( .A(n12069), .B(n12188), .Z(n12072) );
  AND U12004 ( .A(n12321), .B(n12061), .Z(n12188) );
  XOR U12005 ( .A(n12195), .B(n12196), .Z(n12069) );
  ANDN U12006 ( .A(n12197), .B(n12198), .Z(n12196) );
  XNOR U12007 ( .A(n12195), .B(n12199), .Z(n12197) );
  XOR U12008 ( .A(n12078), .B(n12200), .Z(n12073) );
  IV U12009 ( .A(n12077), .Z(n12200) );
  XNOR U12010 ( .A(n12074), .B(n12201), .Z(n12077) );
  XOR U12011 ( .A(n12202), .B(n12203), .Z(n12074) );
  ANDN U12012 ( .A(n12204), .B(n12205), .Z(n12203) );
  XNOR U12013 ( .A(n12202), .B(n12206), .Z(n12204) );
  XNOR U12014 ( .A(n12207), .B(n12208), .Z(n12078) );
  ANDN U12015 ( .A(n12209), .B(n12210), .Z(n12208) );
  XNOR U12016 ( .A(n12207), .B(n12211), .Z(n12209) );
  XOR U12017 ( .A(n12079), .B(n12201), .Z(n12081) );
  AND U12018 ( .A(n11812), .B(n12581), .Z(n12201) );
  XOR U12019 ( .A(n12212), .B(n12213), .Z(n12079) );
  AND U12020 ( .A(n12214), .B(n12215), .Z(n12213) );
  XNOR U12021 ( .A(n12216), .B(n12212), .Z(n12215) );
  XOR U12022 ( .A(n12217), .B(n12181), .Z(n12184) );
  XOR U12023 ( .A(n12218), .B(n12219), .Z(n12181) );
  XNOR U12024 ( .A(n12179), .B(n12182), .Z(n12217) );
  XOR U12025 ( .A(n12220), .B(n12091), .Z(n12179) );
  XOR U12026 ( .A(n12098), .B(n12221), .Z(n12091) );
  IV U12027 ( .A(n12096), .Z(n12221) );
  XNOR U12028 ( .A(n12222), .B(n12095), .Z(n12096) );
  OR U12029 ( .A(n12223), .B(n12224), .Z(n12095) );
  NANDN U12030 ( .B(n6541), .A(n10731), .Z(n12222) );
  XOR U12031 ( .A(n12105), .B(n12225), .Z(n12098) );
  IV U12032 ( .A(n12104), .Z(n12225) );
  XNOR U12033 ( .A(n12101), .B(n12226), .Z(n12104) );
  XOR U12034 ( .A(n12227), .B(n12228), .Z(n12101) );
  NANDN U12035 ( .B(n12229), .A(n12230), .Z(n12227) );
  XOR U12036 ( .A(n12228), .B(n12231), .Z(n12230) );
  XOR U12037 ( .A(n12112), .B(n12232), .Z(n12105) );
  IV U12038 ( .A(n12111), .Z(n12232) );
  XNOR U12039 ( .A(n12108), .B(n12233), .Z(n12111) );
  XOR U12040 ( .A(n12234), .B(n12235), .Z(n12108) );
  ANDN U12041 ( .A(n12236), .B(n12237), .Z(n12235) );
  XNOR U12042 ( .A(n12234), .B(n12238), .Z(n12236) );
  XOR U12043 ( .A(n12119), .B(n12239), .Z(n12112) );
  IV U12044 ( .A(n12118), .Z(n12239) );
  XNOR U12045 ( .A(n12115), .B(n12240), .Z(n12118) );
  XOR U12046 ( .A(n12241), .B(n12242), .Z(n12115) );
  ANDN U12047 ( .A(n12243), .B(n12244), .Z(n12242) );
  XNOR U12048 ( .A(n12241), .B(n12245), .Z(n12243) );
  XOR U12049 ( .A(n12126), .B(n12246), .Z(n12119) );
  IV U12050 ( .A(n12125), .Z(n12246) );
  XNOR U12051 ( .A(n12122), .B(n12247), .Z(n12125) );
  XOR U12052 ( .A(n12248), .B(n12249), .Z(n12122) );
  ANDN U12053 ( .A(n12250), .B(n12251), .Z(n12249) );
  XNOR U12054 ( .A(n12248), .B(n12252), .Z(n12250) );
  XOR U12055 ( .A(n12133), .B(n12253), .Z(n12126) );
  IV U12056 ( .A(n12132), .Z(n12253) );
  XNOR U12057 ( .A(n12129), .B(n12254), .Z(n12132) );
  XOR U12058 ( .A(n12255), .B(n12256), .Z(n12129) );
  ANDN U12059 ( .A(n12257), .B(n12258), .Z(n12256) );
  XNOR U12060 ( .A(n12255), .B(n12259), .Z(n12257) );
  XOR U12061 ( .A(n12139), .B(n12260), .Z(n12133) );
  IV U12062 ( .A(n12138), .Z(n12260) );
  XNOR U12063 ( .A(n12135), .B(n12254), .Z(n12138) );
  AND U12064 ( .A(n12387), .B(n12128), .Z(n12254) );
  XOR U12065 ( .A(n12261), .B(n12262), .Z(n12135) );
  ANDN U12066 ( .A(n12263), .B(n12264), .Z(n12262) );
  XNOR U12067 ( .A(n12261), .B(n12265), .Z(n12263) );
  XOR U12068 ( .A(n12145), .B(n12266), .Z(n12139) );
  IV U12069 ( .A(n12144), .Z(n12266) );
  XNOR U12070 ( .A(n12141), .B(n12247), .Z(n12144) );
  AND U12071 ( .A(n12644), .B(n11869), .Z(n12247) );
  XOR U12072 ( .A(n12267), .B(n12268), .Z(n12141) );
  ANDN U12073 ( .A(n12269), .B(n12270), .Z(n12268) );
  XNOR U12074 ( .A(n12267), .B(n12271), .Z(n12269) );
  XOR U12075 ( .A(n12151), .B(n12272), .Z(n12145) );
  IV U12076 ( .A(n12150), .Z(n12272) );
  XNOR U12077 ( .A(n12147), .B(n12240), .Z(n12150) );
  AND U12078 ( .A(n12880), .B(n11607), .Z(n12240) );
  XOR U12079 ( .A(n12273), .B(n12274), .Z(n12147) );
  ANDN U12080 ( .A(n12275), .B(n12276), .Z(n12274) );
  XNOR U12081 ( .A(n12273), .B(n12277), .Z(n12275) );
  XOR U12082 ( .A(n12157), .B(n12278), .Z(n12151) );
  IV U12083 ( .A(n12156), .Z(n12278) );
  XNOR U12084 ( .A(n12153), .B(n12233), .Z(n12156) );
  AND U12085 ( .A(n13070), .B(n11341), .Z(n12233) );
  XOR U12086 ( .A(n12279), .B(n12280), .Z(n12153) );
  ANDN U12087 ( .A(n12281), .B(n12282), .Z(n12280) );
  XNOR U12088 ( .A(n12279), .B(n12283), .Z(n12281) );
  XOR U12089 ( .A(n12163), .B(n12284), .Z(n12157) );
  IV U12090 ( .A(n12162), .Z(n12284) );
  XNOR U12091 ( .A(n12159), .B(n12226), .Z(n12162) );
  AND U12092 ( .A(n13207), .B(n11049), .Z(n12226) );
  XOR U12093 ( .A(n12285), .B(n12286), .Z(n12159) );
  ANDN U12094 ( .A(n12287), .B(n12288), .Z(n12286) );
  XNOR U12095 ( .A(n12285), .B(n12289), .Z(n12287) );
  XNOR U12096 ( .A(n12168), .B(n12090), .Z(n12163) );
  XNOR U12097 ( .A(n12165), .B(n12290), .Z(n12168) );
  AND U12098 ( .A(n6527), .B(n10731), .Z(n12290) );
  XOR U12099 ( .A(n12291), .B(n12292), .Z(n12165) );
  ANDN U12100 ( .A(n12293), .B(n12294), .Z(n12292) );
  XNOR U12101 ( .A(n12223), .B(n12291), .Z(n12293) );
  XOR U12102 ( .A(n12295), .B(n12090), .Z(n12220) );
  NANDN U12103 ( .B(n6808), .A(n10387), .Z(n12090) );
  XOR U12104 ( .A(n12296), .B(n12297), .Z(n10387) );
  AND U12105 ( .A(n6809), .B(n12298), .Z(n12297) );
  XNOR U12106 ( .A(n12296), .B(n12175), .Z(n12298) );
  XOR U12107 ( .A(n12173), .B(n12296), .Z(n12175) );
  XOR U12108 ( .A(n12299), .B(n12300), .Z(n12173) );
  ANDN U12109 ( .A(n12299), .B(n12301), .Z(n12300) );
  XOR U12110 ( .A(n12302), .B(n7368), .Z(n12296) );
  IV U12111 ( .A(n12177), .Z(n12295) );
  XOR U12112 ( .A(n12303), .B(n12304), .Z(n12177) );
  AND U12113 ( .A(n12305), .B(n12306), .Z(n12304) );
  XNOR U12114 ( .A(n12303), .B(n12307), .Z(n12306) );
  XOR U12115 ( .A(n12308), .B(n12309), .Z(n12182) );
  AND U12116 ( .A(n12310), .B(n12311), .Z(n12309) );
  XOR U12117 ( .A(n12214), .B(n12312), .Z(n12311) );
  XNOR U12118 ( .A(n12308), .B(n12216), .Z(n12312) );
  XOR U12119 ( .A(n12193), .B(n12313), .Z(n12216) );
  IV U12120 ( .A(n12192), .Z(n12313) );
  XNOR U12121 ( .A(n12189), .B(n12314), .Z(n12192) );
  XOR U12122 ( .A(n12315), .B(n12316), .Z(n12189) );
  ANDN U12123 ( .A(n12317), .B(n12318), .Z(n12316) );
  XNOR U12124 ( .A(n12315), .B(n12319), .Z(n12317) );
  XOR U12125 ( .A(n12199), .B(n12320), .Z(n12193) );
  IV U12126 ( .A(n12198), .Z(n12320) );
  XNOR U12127 ( .A(n12195), .B(n12321), .Z(n12198) );
  XOR U12128 ( .A(n12322), .B(n12323), .Z(n12195) );
  ANDN U12129 ( .A(n12324), .B(n12325), .Z(n12323) );
  XNOR U12130 ( .A(n12322), .B(n12326), .Z(n12324) );
  XOR U12131 ( .A(n12206), .B(n12327), .Z(n12199) );
  IV U12132 ( .A(n12205), .Z(n12327) );
  XNOR U12133 ( .A(n12202), .B(n12314), .Z(n12205) );
  AND U12134 ( .A(n12581), .B(n12061), .Z(n12314) );
  XOR U12135 ( .A(n12328), .B(n12329), .Z(n12202) );
  ANDN U12136 ( .A(n12330), .B(n12331), .Z(n12329) );
  XNOR U12137 ( .A(n12328), .B(n12332), .Z(n12330) );
  XOR U12138 ( .A(n12211), .B(n12333), .Z(n12206) );
  IV U12139 ( .A(n12210), .Z(n12333) );
  XNOR U12140 ( .A(n12207), .B(n12334), .Z(n12210) );
  XOR U12141 ( .A(n12335), .B(n12336), .Z(n12207) );
  ANDN U12142 ( .A(n12337), .B(n12338), .Z(n12336) );
  XNOR U12143 ( .A(n12335), .B(n12339), .Z(n12337) );
  XNOR U12144 ( .A(n12340), .B(n12341), .Z(n12211) );
  ANDN U12145 ( .A(n12342), .B(n12343), .Z(n12341) );
  XNOR U12146 ( .A(n12340), .B(n12344), .Z(n12342) );
  XOR U12147 ( .A(n12212), .B(n12334), .Z(n12214) );
  AND U12148 ( .A(n11812), .B(n12827), .Z(n12334) );
  XOR U12149 ( .A(n12345), .B(n12346), .Z(n12212) );
  AND U12150 ( .A(n12347), .B(n12348), .Z(n12346) );
  XNOR U12151 ( .A(n12349), .B(n12345), .Z(n12348) );
  XOR U12152 ( .A(n12350), .B(n12307), .Z(n12310) );
  XOR U12153 ( .A(n12351), .B(n12352), .Z(n12307) );
  XNOR U12154 ( .A(n12305), .B(n12308), .Z(n12350) );
  XOR U12155 ( .A(n12353), .B(n12224), .Z(n12305) );
  XOR U12156 ( .A(n12231), .B(n12354), .Z(n12224) );
  IV U12157 ( .A(n12229), .Z(n12354) );
  XNOR U12158 ( .A(n12355), .B(n12228), .Z(n12229) );
  OR U12159 ( .A(n12356), .B(n12357), .Z(n12228) );
  NANDN U12160 ( .B(n6541), .A(n11049), .Z(n12355) );
  XOR U12161 ( .A(n12238), .B(n12358), .Z(n12231) );
  IV U12162 ( .A(n12237), .Z(n12358) );
  XNOR U12163 ( .A(n12234), .B(n12359), .Z(n12237) );
  XOR U12164 ( .A(n12360), .B(n12361), .Z(n12234) );
  NANDN U12165 ( .B(n12362), .A(n12363), .Z(n12360) );
  XOR U12166 ( .A(n12361), .B(n12364), .Z(n12363) );
  XOR U12167 ( .A(n12245), .B(n12365), .Z(n12238) );
  IV U12168 ( .A(n12244), .Z(n12365) );
  XNOR U12169 ( .A(n12241), .B(n12366), .Z(n12244) );
  XOR U12170 ( .A(n12367), .B(n12368), .Z(n12241) );
  ANDN U12171 ( .A(n12369), .B(n12370), .Z(n12368) );
  XNOR U12172 ( .A(n12367), .B(n12371), .Z(n12369) );
  XOR U12173 ( .A(n12252), .B(n12372), .Z(n12245) );
  IV U12174 ( .A(n12251), .Z(n12372) );
  XNOR U12175 ( .A(n12248), .B(n12373), .Z(n12251) );
  XOR U12176 ( .A(n12374), .B(n12375), .Z(n12248) );
  ANDN U12177 ( .A(n12376), .B(n12377), .Z(n12375) );
  XNOR U12178 ( .A(n12374), .B(n12378), .Z(n12376) );
  XOR U12179 ( .A(n12259), .B(n12379), .Z(n12252) );
  IV U12180 ( .A(n12258), .Z(n12379) );
  XNOR U12181 ( .A(n12255), .B(n12380), .Z(n12258) );
  XOR U12182 ( .A(n12381), .B(n12382), .Z(n12255) );
  ANDN U12183 ( .A(n12383), .B(n12384), .Z(n12382) );
  XNOR U12184 ( .A(n12381), .B(n12385), .Z(n12383) );
  XOR U12185 ( .A(n12265), .B(n12386), .Z(n12259) );
  IV U12186 ( .A(n12264), .Z(n12386) );
  XNOR U12187 ( .A(n12261), .B(n12387), .Z(n12264) );
  XOR U12188 ( .A(n12388), .B(n12389), .Z(n12261) );
  ANDN U12189 ( .A(n12390), .B(n12391), .Z(n12389) );
  XNOR U12190 ( .A(n12388), .B(n12392), .Z(n12390) );
  XOR U12191 ( .A(n12271), .B(n12393), .Z(n12265) );
  IV U12192 ( .A(n12270), .Z(n12393) );
  XNOR U12193 ( .A(n12267), .B(n12380), .Z(n12270) );
  AND U12194 ( .A(n12644), .B(n12128), .Z(n12380) );
  XOR U12195 ( .A(n12394), .B(n12395), .Z(n12267) );
  ANDN U12196 ( .A(n12396), .B(n12397), .Z(n12395) );
  XNOR U12197 ( .A(n12394), .B(n12398), .Z(n12396) );
  XOR U12198 ( .A(n12277), .B(n12399), .Z(n12271) );
  IV U12199 ( .A(n12276), .Z(n12399) );
  XNOR U12200 ( .A(n12273), .B(n12373), .Z(n12276) );
  AND U12201 ( .A(n12880), .B(n11869), .Z(n12373) );
  XOR U12202 ( .A(n12400), .B(n12401), .Z(n12273) );
  ANDN U12203 ( .A(n12402), .B(n12403), .Z(n12401) );
  XNOR U12204 ( .A(n12400), .B(n12404), .Z(n12402) );
  XOR U12205 ( .A(n12283), .B(n12405), .Z(n12277) );
  IV U12206 ( .A(n12282), .Z(n12405) );
  XNOR U12207 ( .A(n12279), .B(n12366), .Z(n12282) );
  AND U12208 ( .A(n13070), .B(n11607), .Z(n12366) );
  XOR U12209 ( .A(n12406), .B(n12407), .Z(n12279) );
  ANDN U12210 ( .A(n12408), .B(n12409), .Z(n12407) );
  XNOR U12211 ( .A(n12406), .B(n12410), .Z(n12408) );
  XOR U12212 ( .A(n12289), .B(n12411), .Z(n12283) );
  IV U12213 ( .A(n12288), .Z(n12411) );
  XNOR U12214 ( .A(n12285), .B(n12359), .Z(n12288) );
  AND U12215 ( .A(n13207), .B(n11341), .Z(n12359) );
  XOR U12216 ( .A(n12412), .B(n12413), .Z(n12285) );
  ANDN U12217 ( .A(n12414), .B(n12415), .Z(n12413) );
  XNOR U12218 ( .A(n12412), .B(n12416), .Z(n12414) );
  XNOR U12219 ( .A(n12294), .B(n12223), .Z(n12289) );
  XNOR U12220 ( .A(n12291), .B(n12417), .Z(n12294) );
  AND U12221 ( .A(n6527), .B(n11049), .Z(n12417) );
  XOR U12222 ( .A(n12418), .B(n12419), .Z(n12291) );
  ANDN U12223 ( .A(n12420), .B(n12421), .Z(n12419) );
  XNOR U12224 ( .A(n12356), .B(n12418), .Z(n12420) );
  XOR U12225 ( .A(n12422), .B(n12223), .Z(n12353) );
  NANDN U12226 ( .B(n6808), .A(n10731), .Z(n12223) );
  XOR U12227 ( .A(n12423), .B(n12424), .Z(n10731) );
  AND U12228 ( .A(n6809), .B(n12425), .Z(n12424) );
  XNOR U12229 ( .A(n12423), .B(n12301), .Z(n12425) );
  XOR U12230 ( .A(n12299), .B(n12423), .Z(n12301) );
  XOR U12231 ( .A(n12426), .B(n12427), .Z(n12299) );
  ANDN U12232 ( .A(n12426), .B(n12428), .Z(n12427) );
  XOR U12233 ( .A(n12429), .B(n7368), .Z(n12423) );
  IV U12234 ( .A(n12303), .Z(n12422) );
  XOR U12235 ( .A(n12430), .B(n12431), .Z(n12303) );
  AND U12236 ( .A(n12432), .B(n12433), .Z(n12431) );
  XNOR U12237 ( .A(n12430), .B(n12434), .Z(n12433) );
  XOR U12238 ( .A(n12435), .B(n12436), .Z(n12308) );
  AND U12239 ( .A(n12437), .B(n12438), .Z(n12436) );
  XOR U12240 ( .A(n12347), .B(n12439), .Z(n12438) );
  XNOR U12241 ( .A(n12435), .B(n12349), .Z(n12439) );
  XOR U12242 ( .A(n12319), .B(n12440), .Z(n12349) );
  IV U12243 ( .A(n12318), .Z(n12440) );
  XNOR U12244 ( .A(n12315), .B(n12441), .Z(n12318) );
  XOR U12245 ( .A(n12442), .B(n12443), .Z(n12315) );
  ANDN U12246 ( .A(n12444), .B(n12445), .Z(n12443) );
  XNOR U12247 ( .A(n12442), .B(n12446), .Z(n12444) );
  XOR U12248 ( .A(n12326), .B(n12447), .Z(n12319) );
  IV U12249 ( .A(n12325), .Z(n12447) );
  XNOR U12250 ( .A(n12322), .B(n12448), .Z(n12325) );
  XOR U12251 ( .A(n12449), .B(n12450), .Z(n12322) );
  ANDN U12252 ( .A(n12451), .B(n12452), .Z(n12450) );
  XNOR U12253 ( .A(n12449), .B(n12453), .Z(n12451) );
  XOR U12254 ( .A(n12332), .B(n12454), .Z(n12326) );
  IV U12255 ( .A(n12331), .Z(n12454) );
  XNOR U12256 ( .A(n12328), .B(n12448), .Z(n12331) );
  AND U12257 ( .A(n12581), .B(n12321), .Z(n12448) );
  XOR U12258 ( .A(n12455), .B(n12456), .Z(n12328) );
  ANDN U12259 ( .A(n12457), .B(n12458), .Z(n12456) );
  XNOR U12260 ( .A(n12455), .B(n12459), .Z(n12457) );
  XOR U12261 ( .A(n12339), .B(n12460), .Z(n12332) );
  IV U12262 ( .A(n12338), .Z(n12460) );
  XNOR U12263 ( .A(n12335), .B(n12441), .Z(n12338) );
  AND U12264 ( .A(n12827), .B(n12061), .Z(n12441) );
  XOR U12265 ( .A(n12461), .B(n12462), .Z(n12335) );
  ANDN U12266 ( .A(n12463), .B(n12464), .Z(n12462) );
  XNOR U12267 ( .A(n12461), .B(n12465), .Z(n12463) );
  XOR U12268 ( .A(n12344), .B(n12466), .Z(n12339) );
  IV U12269 ( .A(n12343), .Z(n12466) );
  XNOR U12270 ( .A(n12340), .B(n12467), .Z(n12343) );
  XOR U12271 ( .A(n12468), .B(n12469), .Z(n12340) );
  ANDN U12272 ( .A(n12470), .B(n12471), .Z(n12469) );
  XNOR U12273 ( .A(n12468), .B(n12472), .Z(n12470) );
  XNOR U12274 ( .A(n12473), .B(n12474), .Z(n12344) );
  ANDN U12275 ( .A(n12475), .B(n12476), .Z(n12474) );
  XNOR U12276 ( .A(n12473), .B(n12477), .Z(n12475) );
  XOR U12277 ( .A(n12345), .B(n12467), .Z(n12347) );
  AND U12278 ( .A(n11812), .B(n13031), .Z(n12467) );
  XOR U12279 ( .A(n12478), .B(n12479), .Z(n12345) );
  AND U12280 ( .A(n12480), .B(n12481), .Z(n12479) );
  XNOR U12281 ( .A(n12482), .B(n12478), .Z(n12481) );
  XOR U12282 ( .A(n12483), .B(n12434), .Z(n12437) );
  XOR U12283 ( .A(n12484), .B(n12485), .Z(n12434) );
  XNOR U12284 ( .A(n12432), .B(n12435), .Z(n12483) );
  XOR U12285 ( .A(n12486), .B(n12357), .Z(n12432) );
  XOR U12286 ( .A(n12364), .B(n12487), .Z(n12357) );
  IV U12287 ( .A(n12362), .Z(n12487) );
  XNOR U12288 ( .A(n12488), .B(n12361), .Z(n12362) );
  OR U12289 ( .A(n12489), .B(n12490), .Z(n12361) );
  NANDN U12290 ( .B(n6541), .A(n11341), .Z(n12488) );
  XOR U12291 ( .A(n12371), .B(n12491), .Z(n12364) );
  IV U12292 ( .A(n12370), .Z(n12491) );
  XNOR U12293 ( .A(n12367), .B(n12492), .Z(n12370) );
  XOR U12294 ( .A(n12493), .B(n12494), .Z(n12367) );
  NANDN U12295 ( .B(n12495), .A(n12496), .Z(n12493) );
  XOR U12296 ( .A(n12494), .B(n12497), .Z(n12496) );
  XOR U12297 ( .A(n12378), .B(n12498), .Z(n12371) );
  IV U12298 ( .A(n12377), .Z(n12498) );
  XNOR U12299 ( .A(n12374), .B(n12499), .Z(n12377) );
  XOR U12300 ( .A(n12500), .B(n12501), .Z(n12374) );
  ANDN U12301 ( .A(n12502), .B(n12503), .Z(n12501) );
  XNOR U12302 ( .A(n12500), .B(n12504), .Z(n12502) );
  XOR U12303 ( .A(n12385), .B(n12505), .Z(n12378) );
  IV U12304 ( .A(n12384), .Z(n12505) );
  XNOR U12305 ( .A(n12381), .B(n12506), .Z(n12384) );
  XOR U12306 ( .A(n12507), .B(n12508), .Z(n12381) );
  ANDN U12307 ( .A(n12509), .B(n12510), .Z(n12508) );
  XNOR U12308 ( .A(n12507), .B(n12511), .Z(n12509) );
  XOR U12309 ( .A(n12392), .B(n12512), .Z(n12385) );
  IV U12310 ( .A(n12391), .Z(n12512) );
  XNOR U12311 ( .A(n12388), .B(n12513), .Z(n12391) );
  XOR U12312 ( .A(n12514), .B(n12515), .Z(n12388) );
  ANDN U12313 ( .A(n12516), .B(n12517), .Z(n12515) );
  XNOR U12314 ( .A(n12514), .B(n12518), .Z(n12516) );
  XOR U12315 ( .A(n12398), .B(n12519), .Z(n12392) );
  IV U12316 ( .A(n12397), .Z(n12519) );
  XNOR U12317 ( .A(n12394), .B(n12513), .Z(n12397) );
  AND U12318 ( .A(n12644), .B(n12387), .Z(n12513) );
  XOR U12319 ( .A(n12520), .B(n12521), .Z(n12394) );
  ANDN U12320 ( .A(n12522), .B(n12523), .Z(n12521) );
  XNOR U12321 ( .A(n12520), .B(n12524), .Z(n12522) );
  XOR U12322 ( .A(n12404), .B(n12525), .Z(n12398) );
  IV U12323 ( .A(n12403), .Z(n12525) );
  XNOR U12324 ( .A(n12400), .B(n12506), .Z(n12403) );
  AND U12325 ( .A(n12880), .B(n12128), .Z(n12506) );
  XOR U12326 ( .A(n12526), .B(n12527), .Z(n12400) );
  ANDN U12327 ( .A(n12528), .B(n12529), .Z(n12527) );
  XNOR U12328 ( .A(n12526), .B(n12530), .Z(n12528) );
  XOR U12329 ( .A(n12410), .B(n12531), .Z(n12404) );
  IV U12330 ( .A(n12409), .Z(n12531) );
  XNOR U12331 ( .A(n12406), .B(n12499), .Z(n12409) );
  AND U12332 ( .A(n13070), .B(n11869), .Z(n12499) );
  XOR U12333 ( .A(n12532), .B(n12533), .Z(n12406) );
  ANDN U12334 ( .A(n12534), .B(n12535), .Z(n12533) );
  XNOR U12335 ( .A(n12532), .B(n12536), .Z(n12534) );
  XOR U12336 ( .A(n12416), .B(n12537), .Z(n12410) );
  IV U12337 ( .A(n12415), .Z(n12537) );
  XNOR U12338 ( .A(n12412), .B(n12492), .Z(n12415) );
  AND U12339 ( .A(n13207), .B(n11607), .Z(n12492) );
  XOR U12340 ( .A(n12538), .B(n12539), .Z(n12412) );
  ANDN U12341 ( .A(n12540), .B(n12541), .Z(n12539) );
  XNOR U12342 ( .A(n12538), .B(n12542), .Z(n12540) );
  XNOR U12343 ( .A(n12421), .B(n12356), .Z(n12416) );
  XNOR U12344 ( .A(n12418), .B(n12543), .Z(n12421) );
  AND U12345 ( .A(n6527), .B(n11341), .Z(n12543) );
  XOR U12346 ( .A(n12544), .B(n12545), .Z(n12418) );
  ANDN U12347 ( .A(n12546), .B(n12547), .Z(n12545) );
  XNOR U12348 ( .A(n12489), .B(n12544), .Z(n12546) );
  XOR U12349 ( .A(n12548), .B(n12356), .Z(n12486) );
  NANDN U12350 ( .B(n6808), .A(n11049), .Z(n12356) );
  XOR U12351 ( .A(n12549), .B(n12550), .Z(n11049) );
  AND U12352 ( .A(n6809), .B(n12551), .Z(n12550) );
  XNOR U12353 ( .A(n12549), .B(n12428), .Z(n12551) );
  XOR U12354 ( .A(n12426), .B(n12549), .Z(n12428) );
  XOR U12355 ( .A(n12552), .B(n12553), .Z(n12426) );
  ANDN U12356 ( .A(n12552), .B(n12554), .Z(n12553) );
  XOR U12357 ( .A(n12555), .B(n7368), .Z(n12549) );
  IV U12358 ( .A(n12430), .Z(n12548) );
  XOR U12359 ( .A(n12556), .B(n12557), .Z(n12430) );
  AND U12360 ( .A(n12558), .B(n12559), .Z(n12557) );
  XNOR U12361 ( .A(n12556), .B(n12560), .Z(n12559) );
  XOR U12362 ( .A(n12561), .B(n12562), .Z(n12435) );
  AND U12363 ( .A(n12563), .B(n12564), .Z(n12562) );
  XOR U12364 ( .A(n12480), .B(n12565), .Z(n12564) );
  XNOR U12365 ( .A(n12561), .B(n12482), .Z(n12565) );
  XOR U12366 ( .A(n12446), .B(n12566), .Z(n12482) );
  IV U12367 ( .A(n12445), .Z(n12566) );
  XNOR U12368 ( .A(n12442), .B(n12567), .Z(n12445) );
  XOR U12369 ( .A(n12568), .B(n12569), .Z(n12442) );
  ANDN U12370 ( .A(n12570), .B(n12571), .Z(n12569) );
  XNOR U12371 ( .A(n12568), .B(n12572), .Z(n12570) );
  XOR U12372 ( .A(n12453), .B(n12573), .Z(n12446) );
  IV U12373 ( .A(n12452), .Z(n12573) );
  XNOR U12374 ( .A(n12449), .B(n12574), .Z(n12452) );
  XOR U12375 ( .A(n12575), .B(n12576), .Z(n12449) );
  ANDN U12376 ( .A(n12577), .B(n12578), .Z(n12576) );
  XNOR U12377 ( .A(n12575), .B(n12579), .Z(n12577) );
  XOR U12378 ( .A(n12459), .B(n12580), .Z(n12453) );
  IV U12379 ( .A(n12458), .Z(n12580) );
  XNOR U12380 ( .A(n12455), .B(n12581), .Z(n12458) );
  XOR U12381 ( .A(n12582), .B(n12583), .Z(n12455) );
  ANDN U12382 ( .A(n12584), .B(n12585), .Z(n12583) );
  XNOR U12383 ( .A(n12582), .B(n12586), .Z(n12584) );
  XOR U12384 ( .A(n12465), .B(n12587), .Z(n12459) );
  IV U12385 ( .A(n12464), .Z(n12587) );
  XNOR U12386 ( .A(n12461), .B(n12574), .Z(n12464) );
  AND U12387 ( .A(n12827), .B(n12321), .Z(n12574) );
  XOR U12388 ( .A(n12588), .B(n12589), .Z(n12461) );
  ANDN U12389 ( .A(n12590), .B(n12591), .Z(n12589) );
  XNOR U12390 ( .A(n12588), .B(n12592), .Z(n12590) );
  XOR U12391 ( .A(n12472), .B(n12593), .Z(n12465) );
  IV U12392 ( .A(n12471), .Z(n12593) );
  XNOR U12393 ( .A(n12468), .B(n12567), .Z(n12471) );
  AND U12394 ( .A(n13031), .B(n12061), .Z(n12567) );
  XOR U12395 ( .A(n12594), .B(n12595), .Z(n12468) );
  ANDN U12396 ( .A(n12596), .B(n12597), .Z(n12595) );
  XNOR U12397 ( .A(n12594), .B(n12598), .Z(n12596) );
  XOR U12398 ( .A(n12477), .B(n12599), .Z(n12472) );
  IV U12399 ( .A(n12476), .Z(n12599) );
  XNOR U12400 ( .A(n12473), .B(n12600), .Z(n12476) );
  XOR U12401 ( .A(n12601), .B(n12602), .Z(n12473) );
  ANDN U12402 ( .A(n12603), .B(n12604), .Z(n12602) );
  XOR U12403 ( .A(n12601), .B(n12605), .Z(n12603) );
  XNOR U12404 ( .A(n12606), .B(n12607), .Z(n12477) );
  ANDN U12405 ( .A(n12606), .B(n12608), .Z(n12607) );
  XOR U12406 ( .A(n12478), .B(n12600), .Z(n12480) );
  AND U12407 ( .A(n11812), .B(n13181), .Z(n12600) );
  XOR U12408 ( .A(n12609), .B(n12610), .Z(n12478) );
  NAND U12409 ( .A(n12611), .B(n12612), .Z(n12609) );
  XOR U12410 ( .A(n12610), .B(n12613), .Z(n12611) );
  XOR U12411 ( .A(n12614), .B(n12560), .Z(n12563) );
  XOR U12412 ( .A(n12615), .B(n12616), .Z(n12560) );
  XNOR U12413 ( .A(n12558), .B(n12561), .Z(n12614) );
  XOR U12414 ( .A(n12617), .B(n12490), .Z(n12558) );
  XOR U12415 ( .A(n12497), .B(n12618), .Z(n12490) );
  IV U12416 ( .A(n12495), .Z(n12618) );
  XNOR U12417 ( .A(n12619), .B(n12494), .Z(n12495) );
  OR U12418 ( .A(n12620), .B(n12621), .Z(n12494) );
  NANDN U12419 ( .B(n6541), .A(n11607), .Z(n12619) );
  XOR U12420 ( .A(n12504), .B(n12622), .Z(n12497) );
  IV U12421 ( .A(n12503), .Z(n12622) );
  XNOR U12422 ( .A(n12500), .B(n12623), .Z(n12503) );
  XOR U12423 ( .A(n12624), .B(n12625), .Z(n12500) );
  NANDN U12424 ( .B(n12626), .A(n12627), .Z(n12624) );
  XOR U12425 ( .A(n12625), .B(n12628), .Z(n12627) );
  XOR U12426 ( .A(n12511), .B(n12629), .Z(n12504) );
  IV U12427 ( .A(n12510), .Z(n12629) );
  XNOR U12428 ( .A(n12507), .B(n12630), .Z(n12510) );
  XOR U12429 ( .A(n12631), .B(n12632), .Z(n12507) );
  ANDN U12430 ( .A(n12633), .B(n12634), .Z(n12632) );
  XNOR U12431 ( .A(n12631), .B(n12635), .Z(n12633) );
  XOR U12432 ( .A(n12518), .B(n12636), .Z(n12511) );
  IV U12433 ( .A(n12517), .Z(n12636) );
  XNOR U12434 ( .A(n12514), .B(n12637), .Z(n12517) );
  XOR U12435 ( .A(n12638), .B(n12639), .Z(n12514) );
  ANDN U12436 ( .A(n12640), .B(n12641), .Z(n12639) );
  XNOR U12437 ( .A(n12638), .B(n12642), .Z(n12640) );
  XOR U12438 ( .A(n12524), .B(n12643), .Z(n12518) );
  IV U12439 ( .A(n12523), .Z(n12643) );
  XNOR U12440 ( .A(n12520), .B(n12644), .Z(n12523) );
  XOR U12441 ( .A(n12645), .B(n12646), .Z(n12520) );
  ANDN U12442 ( .A(n12647), .B(n12648), .Z(n12646) );
  XNOR U12443 ( .A(n12645), .B(n12649), .Z(n12647) );
  XOR U12444 ( .A(n12530), .B(n12650), .Z(n12524) );
  IV U12445 ( .A(n12529), .Z(n12650) );
  XNOR U12446 ( .A(n12526), .B(n12637), .Z(n12529) );
  AND U12447 ( .A(n12880), .B(n12387), .Z(n12637) );
  XOR U12448 ( .A(n12651), .B(n12652), .Z(n12526) );
  ANDN U12449 ( .A(n12653), .B(n12654), .Z(n12652) );
  XNOR U12450 ( .A(n12651), .B(n12655), .Z(n12653) );
  XOR U12451 ( .A(n12536), .B(n12656), .Z(n12530) );
  IV U12452 ( .A(n12535), .Z(n12656) );
  XNOR U12453 ( .A(n12532), .B(n12630), .Z(n12535) );
  AND U12454 ( .A(n13070), .B(n12128), .Z(n12630) );
  XOR U12455 ( .A(n12657), .B(n12658), .Z(n12532) );
  ANDN U12456 ( .A(n12659), .B(n12660), .Z(n12658) );
  XNOR U12457 ( .A(n12657), .B(n12661), .Z(n12659) );
  XOR U12458 ( .A(n12542), .B(n12662), .Z(n12536) );
  IV U12459 ( .A(n12541), .Z(n12662) );
  XNOR U12460 ( .A(n12538), .B(n12623), .Z(n12541) );
  AND U12461 ( .A(n13207), .B(n11869), .Z(n12623) );
  XOR U12462 ( .A(n12663), .B(n12664), .Z(n12538) );
  ANDN U12463 ( .A(n12665), .B(n12666), .Z(n12664) );
  XNOR U12464 ( .A(n12663), .B(n12667), .Z(n12665) );
  XNOR U12465 ( .A(n12547), .B(n12489), .Z(n12542) );
  XNOR U12466 ( .A(n12544), .B(n12668), .Z(n12547) );
  AND U12467 ( .A(n6527), .B(n11607), .Z(n12668) );
  XOR U12468 ( .A(n12669), .B(n12670), .Z(n12544) );
  ANDN U12469 ( .A(n12671), .B(n12672), .Z(n12670) );
  XNOR U12470 ( .A(n12620), .B(n12669), .Z(n12671) );
  XOR U12471 ( .A(n12673), .B(n12489), .Z(n12617) );
  NANDN U12472 ( .B(n6808), .A(n11341), .Z(n12489) );
  XOR U12473 ( .A(n12674), .B(n12675), .Z(n11341) );
  AND U12474 ( .A(n6809), .B(n12676), .Z(n12675) );
  XNOR U12475 ( .A(n12674), .B(n12554), .Z(n12676) );
  XOR U12476 ( .A(n12552), .B(n12674), .Z(n12554) );
  XOR U12477 ( .A(n12677), .B(n12678), .Z(n12552) );
  ANDN U12478 ( .A(n12677), .B(n12679), .Z(n12678) );
  XOR U12479 ( .A(n12680), .B(n7368), .Z(n12674) );
  IV U12480 ( .A(n12556), .Z(n12673) );
  XOR U12481 ( .A(n12681), .B(n12682), .Z(n12556) );
  AND U12482 ( .A(n12683), .B(n12684), .Z(n12682) );
  XNOR U12483 ( .A(n12681), .B(n12685), .Z(n12684) );
  XOR U12484 ( .A(n12686), .B(n12687), .Z(n12561) );
  AND U12485 ( .A(n12688), .B(n12689), .Z(n12687) );
  XOR U12486 ( .A(n12612), .B(n12690), .Z(n12689) );
  XNOR U12487 ( .A(n12686), .B(n12613), .Z(n12690) );
  XOR U12488 ( .A(n12572), .B(n12691), .Z(n12613) );
  IV U12489 ( .A(n12571), .Z(n12691) );
  XNOR U12490 ( .A(n12568), .B(n12692), .Z(n12571) );
  XOR U12491 ( .A(n12693), .B(n12694), .Z(n12568) );
  NANDN U12492 ( .B(n12695), .A(n12696), .Z(n12693) );
  XOR U12493 ( .A(n12694), .B(n12697), .Z(n12696) );
  XOR U12494 ( .A(n12579), .B(n12698), .Z(n12572) );
  IV U12495 ( .A(n12578), .Z(n12698) );
  XNOR U12496 ( .A(n12575), .B(n12699), .Z(n12578) );
  XOR U12497 ( .A(n12700), .B(n12701), .Z(n12575) );
  ANDN U12498 ( .A(n12702), .B(n12703), .Z(n12701) );
  XNOR U12499 ( .A(n12700), .B(n12704), .Z(n12702) );
  XOR U12500 ( .A(n12586), .B(n12705), .Z(n12579) );
  IV U12501 ( .A(n12585), .Z(n12705) );
  XNOR U12502 ( .A(n12582), .B(n12706), .Z(n12585) );
  XOR U12503 ( .A(n12707), .B(n12708), .Z(n12582) );
  ANDN U12504 ( .A(n12709), .B(n12710), .Z(n12708) );
  XNOR U12505 ( .A(n12707), .B(n12711), .Z(n12709) );
  XOR U12506 ( .A(n12592), .B(n12712), .Z(n12586) );
  IV U12507 ( .A(n12591), .Z(n12712) );
  XNOR U12508 ( .A(n12588), .B(n12706), .Z(n12591) );
  AND U12509 ( .A(n12827), .B(n12581), .Z(n12706) );
  XOR U12510 ( .A(n12713), .B(n12714), .Z(n12588) );
  ANDN U12511 ( .A(n12715), .B(n12716), .Z(n12714) );
  XNOR U12512 ( .A(n12713), .B(n12717), .Z(n12715) );
  XOR U12513 ( .A(n12598), .B(n12718), .Z(n12592) );
  IV U12514 ( .A(n12597), .Z(n12718) );
  XNOR U12515 ( .A(n12594), .B(n12699), .Z(n12597) );
  AND U12516 ( .A(n13031), .B(n12321), .Z(n12699) );
  XOR U12517 ( .A(n12719), .B(n12720), .Z(n12594) );
  ANDN U12518 ( .A(n12721), .B(n12722), .Z(n12720) );
  XNOR U12519 ( .A(n12719), .B(n12723), .Z(n12721) );
  XOR U12520 ( .A(n12605), .B(n12604), .Z(n12598) );
  XNOR U12521 ( .A(n12601), .B(n12692), .Z(n12604) );
  AND U12522 ( .A(n13181), .B(n12061), .Z(n12692) );
  XOR U12523 ( .A(n12724), .B(n12725), .Z(n12601) );
  ANDN U12524 ( .A(n12726), .B(n12727), .Z(n12725) );
  XNOR U12525 ( .A(n12724), .B(n12728), .Z(n12726) );
  IV U12526 ( .A(n12608), .Z(n12605) );
  XNOR U12527 ( .A(n12606), .B(n12729), .Z(n12608) );
  AND U12528 ( .A(n11812), .B(n12730), .Z(n12729) );
  XOR U12529 ( .A(n12731), .B(n12732), .Z(n12606) );
  ANDN U12530 ( .A(n12733), .B(n12734), .Z(n12732) );
  XNOR U12531 ( .A(n12735), .B(n12731), .Z(n12733) );
  XOR U12532 ( .A(n12736), .B(n12610), .Z(n12612) );
  OR U12533 ( .A(n12735), .B(n12737), .Z(n12610) );
  NAND U12534 ( .A(n12730), .B(n11812), .Z(n12736) );
  XOR U12535 ( .A(n12738), .B(n12685), .Z(n12688) );
  XOR U12536 ( .A(n12739), .B(n12740), .Z(n12685) );
  XNOR U12537 ( .A(n12683), .B(n12686), .Z(n12738) );
  XOR U12538 ( .A(n12741), .B(n12621), .Z(n12683) );
  XOR U12539 ( .A(n12628), .B(n12742), .Z(n12621) );
  IV U12540 ( .A(n12626), .Z(n12742) );
  XNOR U12541 ( .A(n12743), .B(n12625), .Z(n12626) );
  OR U12542 ( .A(n12744), .B(n12745), .Z(n12625) );
  NANDN U12543 ( .B(n6541), .A(n11869), .Z(n12743) );
  XOR U12544 ( .A(n12635), .B(n12746), .Z(n12628) );
  IV U12545 ( .A(n12634), .Z(n12746) );
  XNOR U12546 ( .A(n12631), .B(n12747), .Z(n12634) );
  XOR U12547 ( .A(n12748), .B(n12749), .Z(n12631) );
  NANDN U12548 ( .B(n12750), .A(n12751), .Z(n12748) );
  XOR U12549 ( .A(n12749), .B(n12752), .Z(n12751) );
  XOR U12550 ( .A(n12642), .B(n12753), .Z(n12635) );
  IV U12551 ( .A(n12641), .Z(n12753) );
  XNOR U12552 ( .A(n12638), .B(n12754), .Z(n12641) );
  XOR U12553 ( .A(n12755), .B(n12756), .Z(n12638) );
  ANDN U12554 ( .A(n12757), .B(n12758), .Z(n12756) );
  XNOR U12555 ( .A(n12755), .B(n12759), .Z(n12757) );
  XOR U12556 ( .A(n12649), .B(n12760), .Z(n12642) );
  IV U12557 ( .A(n12648), .Z(n12760) );
  XNOR U12558 ( .A(n12645), .B(n12761), .Z(n12648) );
  XOR U12559 ( .A(n12762), .B(n12763), .Z(n12645) );
  ANDN U12560 ( .A(n12764), .B(n12765), .Z(n12763) );
  XNOR U12561 ( .A(n12762), .B(n12766), .Z(n12764) );
  XOR U12562 ( .A(n12655), .B(n12767), .Z(n12649) );
  IV U12563 ( .A(n12654), .Z(n12767) );
  XNOR U12564 ( .A(n12651), .B(n12761), .Z(n12654) );
  AND U12565 ( .A(n12880), .B(n12644), .Z(n12761) );
  XOR U12566 ( .A(n12768), .B(n12769), .Z(n12651) );
  ANDN U12567 ( .A(n12770), .B(n12771), .Z(n12769) );
  XNOR U12568 ( .A(n12768), .B(n12772), .Z(n12770) );
  XOR U12569 ( .A(n12661), .B(n12773), .Z(n12655) );
  IV U12570 ( .A(n12660), .Z(n12773) );
  XNOR U12571 ( .A(n12657), .B(n12754), .Z(n12660) );
  AND U12572 ( .A(n13070), .B(n12387), .Z(n12754) );
  XOR U12573 ( .A(n12774), .B(n12775), .Z(n12657) );
  ANDN U12574 ( .A(n12776), .B(n12777), .Z(n12775) );
  XNOR U12575 ( .A(n12774), .B(n12778), .Z(n12776) );
  XOR U12576 ( .A(n12667), .B(n12779), .Z(n12661) );
  IV U12577 ( .A(n12666), .Z(n12779) );
  XNOR U12578 ( .A(n12663), .B(n12747), .Z(n12666) );
  AND U12579 ( .A(n13207), .B(n12128), .Z(n12747) );
  XOR U12580 ( .A(n12780), .B(n12781), .Z(n12663) );
  ANDN U12581 ( .A(n12782), .B(n12783), .Z(n12781) );
  XNOR U12582 ( .A(n12780), .B(n12784), .Z(n12782) );
  XNOR U12583 ( .A(n12672), .B(n12620), .Z(n12667) );
  XNOR U12584 ( .A(n12669), .B(n12785), .Z(n12672) );
  AND U12585 ( .A(n6527), .B(n11869), .Z(n12785) );
  XOR U12586 ( .A(n12786), .B(n12787), .Z(n12669) );
  ANDN U12587 ( .A(n12788), .B(n12789), .Z(n12787) );
  XNOR U12588 ( .A(n12744), .B(n12786), .Z(n12788) );
  XOR U12589 ( .A(n12790), .B(n12620), .Z(n12741) );
  NANDN U12590 ( .B(n6808), .A(n11607), .Z(n12620) );
  XOR U12591 ( .A(n12791), .B(n12792), .Z(n11607) );
  AND U12592 ( .A(n6809), .B(n12793), .Z(n12792) );
  XNOR U12593 ( .A(n12791), .B(n12679), .Z(n12793) );
  XOR U12594 ( .A(n12677), .B(n12791), .Z(n12679) );
  XOR U12595 ( .A(n12794), .B(n12795), .Z(n12677) );
  ANDN U12596 ( .A(n12794), .B(n12796), .Z(n12795) );
  XOR U12597 ( .A(n12797), .B(n7368), .Z(n12791) );
  IV U12598 ( .A(n12681), .Z(n12790) );
  XOR U12599 ( .A(n12798), .B(n12799), .Z(n12681) );
  AND U12600 ( .A(n12800), .B(n12801), .Z(n12799) );
  XNOR U12601 ( .A(n12798), .B(n12802), .Z(n12801) );
  XOR U12602 ( .A(n12803), .B(n12804), .Z(n12686) );
  AND U12603 ( .A(n12805), .B(n12806), .Z(n12804) );
  XNOR U12604 ( .A(n12737), .B(n12807), .Z(n12806) );
  XNOR U12605 ( .A(n12735), .B(n12803), .Z(n12807) );
  XOR U12606 ( .A(n12697), .B(n12808), .Z(n12737) );
  IV U12607 ( .A(n12695), .Z(n12808) );
  XNOR U12608 ( .A(n12809), .B(n12694), .Z(n12695) );
  OR U12609 ( .A(n12810), .B(n12811), .Z(n12694) );
  NAND U12610 ( .A(n12730), .B(n12061), .Z(n12809) );
  XOR U12611 ( .A(n12704), .B(n12812), .Z(n12697) );
  IV U12612 ( .A(n12703), .Z(n12812) );
  XNOR U12613 ( .A(n12700), .B(n12813), .Z(n12703) );
  XOR U12614 ( .A(n12814), .B(n12815), .Z(n12700) );
  NANDN U12615 ( .B(n12816), .A(n12817), .Z(n12814) );
  XOR U12616 ( .A(n12815), .B(n12818), .Z(n12817) );
  XOR U12617 ( .A(n12711), .B(n12819), .Z(n12704) );
  IV U12618 ( .A(n12710), .Z(n12819) );
  XNOR U12619 ( .A(n12707), .B(n12820), .Z(n12710) );
  XOR U12620 ( .A(n12821), .B(n12822), .Z(n12707) );
  ANDN U12621 ( .A(n12823), .B(n12824), .Z(n12822) );
  XNOR U12622 ( .A(n12821), .B(n12825), .Z(n12823) );
  XOR U12623 ( .A(n12717), .B(n12826), .Z(n12711) );
  IV U12624 ( .A(n12716), .Z(n12826) );
  XNOR U12625 ( .A(n12713), .B(n12827), .Z(n12716) );
  XOR U12626 ( .A(n12828), .B(n12829), .Z(n12713) );
  ANDN U12627 ( .A(n12830), .B(n12831), .Z(n12829) );
  XNOR U12628 ( .A(n12828), .B(n12832), .Z(n12830) );
  XOR U12629 ( .A(n12723), .B(n12833), .Z(n12717) );
  IV U12630 ( .A(n12722), .Z(n12833) );
  XNOR U12631 ( .A(n12719), .B(n12820), .Z(n12722) );
  AND U12632 ( .A(n13031), .B(n12581), .Z(n12820) );
  XOR U12633 ( .A(n12834), .B(n12835), .Z(n12719) );
  ANDN U12634 ( .A(n12836), .B(n12837), .Z(n12835) );
  XNOR U12635 ( .A(n12834), .B(n12838), .Z(n12836) );
  XOR U12636 ( .A(n12728), .B(n12839), .Z(n12723) );
  IV U12637 ( .A(n12727), .Z(n12839) );
  XNOR U12638 ( .A(n12724), .B(n12813), .Z(n12727) );
  AND U12639 ( .A(n13181), .B(n12321), .Z(n12813) );
  XOR U12640 ( .A(n12840), .B(n12841), .Z(n12724) );
  ANDN U12641 ( .A(n12842), .B(n12843), .Z(n12841) );
  XNOR U12642 ( .A(n12840), .B(n12844), .Z(n12842) );
  XNOR U12643 ( .A(n12734), .B(n12735), .Z(n12728) );
  NANDN U12644 ( .B(n12845), .A(n11812), .Z(n12735) );
  XNOR U12645 ( .A(n12846), .B(e_input[8]), .Z(n11812) );
  NANDN U12646 ( .B(n12847), .A(n12848), .Z(n12846) );
  XNOR U12647 ( .A(n12849), .B(n12850), .Z(n12848) );
  ANDN U12648 ( .A(n12850), .B(n12851), .Z(n12849) );
  XNOR U12649 ( .A(n12731), .B(n12852), .Z(n12734) );
  AND U12650 ( .A(n12730), .B(n12061), .Z(n12852) );
  XOR U12651 ( .A(n12853), .B(n12854), .Z(n12731) );
  ANDN U12652 ( .A(n12855), .B(n12856), .Z(n12854) );
  XNOR U12653 ( .A(n12810), .B(n12853), .Z(n12855) );
  XOR U12654 ( .A(n12857), .B(n12802), .Z(n12805) );
  XOR U12655 ( .A(n12858), .B(n12859), .Z(n12802) );
  XNOR U12656 ( .A(n12800), .B(n12803), .Z(n12857) );
  XOR U12657 ( .A(n12860), .B(n12745), .Z(n12800) );
  XOR U12658 ( .A(n12752), .B(n12861), .Z(n12745) );
  IV U12659 ( .A(n12750), .Z(n12861) );
  XNOR U12660 ( .A(n12862), .B(n12749), .Z(n12750) );
  OR U12661 ( .A(n12863), .B(n12864), .Z(n12749) );
  NANDN U12662 ( .B(n6541), .A(n12128), .Z(n12862) );
  XOR U12663 ( .A(n12759), .B(n12865), .Z(n12752) );
  IV U12664 ( .A(n12758), .Z(n12865) );
  XNOR U12665 ( .A(n12755), .B(n12866), .Z(n12758) );
  XOR U12666 ( .A(n12867), .B(n12868), .Z(n12755) );
  NANDN U12667 ( .B(n12869), .A(n12870), .Z(n12867) );
  XOR U12668 ( .A(n12868), .B(n12871), .Z(n12870) );
  XOR U12669 ( .A(n12766), .B(n12872), .Z(n12759) );
  IV U12670 ( .A(n12765), .Z(n12872) );
  XNOR U12671 ( .A(n12762), .B(n12873), .Z(n12765) );
  XOR U12672 ( .A(n12874), .B(n12875), .Z(n12762) );
  ANDN U12673 ( .A(n12876), .B(n12877), .Z(n12875) );
  XNOR U12674 ( .A(n12874), .B(n12878), .Z(n12876) );
  XOR U12675 ( .A(n12772), .B(n12879), .Z(n12766) );
  IV U12676 ( .A(n12771), .Z(n12879) );
  XNOR U12677 ( .A(n12768), .B(n12880), .Z(n12771) );
  XOR U12678 ( .A(n12881), .B(n12882), .Z(n12768) );
  ANDN U12679 ( .A(n12883), .B(n12884), .Z(n12882) );
  XNOR U12680 ( .A(n12881), .B(n12885), .Z(n12883) );
  XOR U12681 ( .A(n12778), .B(n12886), .Z(n12772) );
  IV U12682 ( .A(n12777), .Z(n12886) );
  XNOR U12683 ( .A(n12774), .B(n12873), .Z(n12777) );
  AND U12684 ( .A(n13070), .B(n12644), .Z(n12873) );
  XOR U12685 ( .A(n12887), .B(n12888), .Z(n12774) );
  ANDN U12686 ( .A(n12889), .B(n12890), .Z(n12888) );
  XNOR U12687 ( .A(n12887), .B(n12891), .Z(n12889) );
  XOR U12688 ( .A(n12784), .B(n12892), .Z(n12778) );
  IV U12689 ( .A(n12783), .Z(n12892) );
  XNOR U12690 ( .A(n12780), .B(n12866), .Z(n12783) );
  AND U12691 ( .A(n13207), .B(n12387), .Z(n12866) );
  XOR U12692 ( .A(n12893), .B(n12894), .Z(n12780) );
  ANDN U12693 ( .A(n12895), .B(n12896), .Z(n12894) );
  XNOR U12694 ( .A(n12893), .B(n12897), .Z(n12895) );
  XNOR U12695 ( .A(n12789), .B(n12744), .Z(n12784) );
  XNOR U12696 ( .A(n12786), .B(n12898), .Z(n12789) );
  AND U12697 ( .A(n6527), .B(n12128), .Z(n12898) );
  XOR U12698 ( .A(n12899), .B(n12900), .Z(n12786) );
  ANDN U12699 ( .A(n12901), .B(n12902), .Z(n12900) );
  XNOR U12700 ( .A(n12863), .B(n12899), .Z(n12901) );
  XOR U12701 ( .A(n12903), .B(n12744), .Z(n12860) );
  NANDN U12702 ( .B(n6808), .A(n11869), .Z(n12744) );
  XOR U12703 ( .A(n12904), .B(n12905), .Z(n11869) );
  AND U12704 ( .A(n6809), .B(n12906), .Z(n12905) );
  XNOR U12705 ( .A(n12904), .B(n12796), .Z(n12906) );
  XOR U12706 ( .A(n12794), .B(n12904), .Z(n12796) );
  XOR U12707 ( .A(n12907), .B(n12908), .Z(n12794) );
  ANDN U12708 ( .A(n12907), .B(n12909), .Z(n12908) );
  XOR U12709 ( .A(n12910), .B(n7368), .Z(n12904) );
  IV U12710 ( .A(n12798), .Z(n12903) );
  XOR U12711 ( .A(n12911), .B(n12912), .Z(n12798) );
  AND U12712 ( .A(n12913), .B(n12914), .Z(n12912) );
  XNOR U12713 ( .A(n12911), .B(n12915), .Z(n12914) );
  XOR U12714 ( .A(n12916), .B(n12917), .Z(n12803) );
  AND U12715 ( .A(n12918), .B(n12919), .Z(n12917) );
  XNOR U12716 ( .A(n12811), .B(n12920), .Z(n12919) );
  XNOR U12717 ( .A(n12810), .B(n12916), .Z(n12920) );
  XOR U12718 ( .A(n12818), .B(n12921), .Z(n12811) );
  IV U12719 ( .A(n12816), .Z(n12921) );
  XNOR U12720 ( .A(n12922), .B(n12815), .Z(n12816) );
  OR U12721 ( .A(n12923), .B(n12924), .Z(n12815) );
  NAND U12722 ( .A(n12730), .B(n12321), .Z(n12922) );
  XOR U12723 ( .A(n12825), .B(n12925), .Z(n12818) );
  IV U12724 ( .A(n12824), .Z(n12925) );
  XNOR U12725 ( .A(n12821), .B(n12926), .Z(n12824) );
  XOR U12726 ( .A(n12927), .B(n12928), .Z(n12821) );
  NANDN U12727 ( .B(n12929), .A(n12930), .Z(n12927) );
  XOR U12728 ( .A(n12928), .B(n12931), .Z(n12930) );
  XOR U12729 ( .A(n12832), .B(n12932), .Z(n12825) );
  IV U12730 ( .A(n12831), .Z(n12932) );
  XNOR U12731 ( .A(n12828), .B(n12933), .Z(n12831) );
  XOR U12732 ( .A(n12934), .B(n12935), .Z(n12828) );
  ANDN U12733 ( .A(n12936), .B(n12937), .Z(n12935) );
  XNOR U12734 ( .A(n12934), .B(n12938), .Z(n12936) );
  XOR U12735 ( .A(n12838), .B(n12939), .Z(n12832) );
  IV U12736 ( .A(n12837), .Z(n12939) );
  XNOR U12737 ( .A(n12834), .B(n12933), .Z(n12837) );
  AND U12738 ( .A(n13031), .B(n12827), .Z(n12933) );
  XOR U12739 ( .A(n12940), .B(n12941), .Z(n12834) );
  ANDN U12740 ( .A(n12942), .B(n12943), .Z(n12941) );
  XNOR U12741 ( .A(n12940), .B(n12944), .Z(n12942) );
  XOR U12742 ( .A(n12844), .B(n12945), .Z(n12838) );
  IV U12743 ( .A(n12843), .Z(n12945) );
  XNOR U12744 ( .A(n12840), .B(n12926), .Z(n12843) );
  AND U12745 ( .A(n13181), .B(n12581), .Z(n12926) );
  XOR U12746 ( .A(n12946), .B(n12947), .Z(n12840) );
  ANDN U12747 ( .A(n12948), .B(n12949), .Z(n12947) );
  XNOR U12748 ( .A(n12946), .B(n12950), .Z(n12948) );
  XNOR U12749 ( .A(n12856), .B(n12810), .Z(n12844) );
  NANDN U12750 ( .B(n12845), .A(n12061), .Z(n12810) );
  XNOR U12751 ( .A(n12951), .B(e_input[7]), .Z(n12061) );
  NANDN U12752 ( .B(n12847), .A(n12952), .Z(n12951) );
  XOR U12753 ( .A(n12953), .B(n12851), .Z(n12952) );
  XNOR U12754 ( .A(n12850), .B(n12953), .Z(n12851) );
  XOR U12755 ( .A(n12954), .B(n12955), .Z(n12850) );
  ANDN U12756 ( .A(n12954), .B(n12956), .Z(n12955) );
  IV U12757 ( .A(e_input[7]), .Z(n12953) );
  XNOR U12758 ( .A(n12853), .B(n12957), .Z(n12856) );
  AND U12759 ( .A(n12730), .B(n12321), .Z(n12957) );
  XOR U12760 ( .A(n12958), .B(n12959), .Z(n12853) );
  ANDN U12761 ( .A(n12960), .B(n12961), .Z(n12959) );
  XNOR U12762 ( .A(n12923), .B(n12958), .Z(n12960) );
  XOR U12763 ( .A(n12962), .B(n12915), .Z(n12918) );
  XOR U12764 ( .A(n12963), .B(n12964), .Z(n12915) );
  XNOR U12765 ( .A(n12913), .B(n12916), .Z(n12962) );
  XOR U12766 ( .A(n12965), .B(n12864), .Z(n12913) );
  XOR U12767 ( .A(n12871), .B(n12966), .Z(n12864) );
  IV U12768 ( .A(n12869), .Z(n12966) );
  XNOR U12769 ( .A(n12967), .B(n12868), .Z(n12869) );
  OR U12770 ( .A(n12968), .B(n12969), .Z(n12868) );
  NANDN U12771 ( .B(n6541), .A(n12387), .Z(n12967) );
  XOR U12772 ( .A(n12878), .B(n12970), .Z(n12871) );
  IV U12773 ( .A(n12877), .Z(n12970) );
  XNOR U12774 ( .A(n12874), .B(n12971), .Z(n12877) );
  XOR U12775 ( .A(n12972), .B(n12973), .Z(n12874) );
  NANDN U12776 ( .B(n12974), .A(n12975), .Z(n12972) );
  XOR U12777 ( .A(n12973), .B(n12976), .Z(n12975) );
  XOR U12778 ( .A(n12885), .B(n12977), .Z(n12878) );
  IV U12779 ( .A(n12884), .Z(n12977) );
  XNOR U12780 ( .A(n12881), .B(n12978), .Z(n12884) );
  XOR U12781 ( .A(n12979), .B(n12980), .Z(n12881) );
  ANDN U12782 ( .A(n12981), .B(n12982), .Z(n12980) );
  XNOR U12783 ( .A(n12979), .B(n12983), .Z(n12981) );
  XOR U12784 ( .A(n12891), .B(n12984), .Z(n12885) );
  IV U12785 ( .A(n12890), .Z(n12984) );
  XNOR U12786 ( .A(n12887), .B(n12978), .Z(n12890) );
  AND U12787 ( .A(n13070), .B(n12880), .Z(n12978) );
  XOR U12788 ( .A(n12985), .B(n12986), .Z(n12887) );
  ANDN U12789 ( .A(n12987), .B(n12988), .Z(n12986) );
  XNOR U12790 ( .A(n12985), .B(n12989), .Z(n12987) );
  XOR U12791 ( .A(n12897), .B(n12990), .Z(n12891) );
  IV U12792 ( .A(n12896), .Z(n12990) );
  XNOR U12793 ( .A(n12893), .B(n12971), .Z(n12896) );
  AND U12794 ( .A(n13207), .B(n12644), .Z(n12971) );
  XOR U12795 ( .A(n12991), .B(n12992), .Z(n12893) );
  ANDN U12796 ( .A(n12993), .B(n12994), .Z(n12992) );
  XNOR U12797 ( .A(n12991), .B(n12995), .Z(n12993) );
  XNOR U12798 ( .A(n12902), .B(n12863), .Z(n12897) );
  XNOR U12799 ( .A(n12899), .B(n12996), .Z(n12902) );
  AND U12800 ( .A(n6527), .B(n12387), .Z(n12996) );
  XOR U12801 ( .A(n12997), .B(n12998), .Z(n12899) );
  ANDN U12802 ( .A(n12999), .B(n13000), .Z(n12998) );
  XNOR U12803 ( .A(n12968), .B(n12997), .Z(n12999) );
  XOR U12804 ( .A(n13001), .B(n12863), .Z(n12965) );
  NANDN U12805 ( .B(n6808), .A(n12128), .Z(n12863) );
  XOR U12806 ( .A(n13002), .B(n13003), .Z(n12128) );
  AND U12807 ( .A(n6809), .B(n13004), .Z(n13003) );
  XNOR U12808 ( .A(n13002), .B(n12909), .Z(n13004) );
  XOR U12809 ( .A(n12907), .B(n13002), .Z(n12909) );
  XOR U12810 ( .A(n13005), .B(n13006), .Z(n12907) );
  ANDN U12811 ( .A(n13005), .B(n13007), .Z(n13006) );
  XOR U12812 ( .A(n13008), .B(n7368), .Z(n13002) );
  IV U12813 ( .A(n12911), .Z(n13001) );
  XOR U12814 ( .A(n13009), .B(n13010), .Z(n12911) );
  AND U12815 ( .A(n13011), .B(n13012), .Z(n13010) );
  XNOR U12816 ( .A(n13009), .B(n13013), .Z(n13012) );
  XOR U12817 ( .A(n13014), .B(n13015), .Z(n12916) );
  AND U12818 ( .A(n13016), .B(n13017), .Z(n13015) );
  XNOR U12819 ( .A(n12924), .B(n13018), .Z(n13017) );
  XNOR U12820 ( .A(n12923), .B(n13014), .Z(n13018) );
  XOR U12821 ( .A(n12931), .B(n13019), .Z(n12924) );
  IV U12822 ( .A(n12929), .Z(n13019) );
  XNOR U12823 ( .A(n13020), .B(n12928), .Z(n12929) );
  OR U12824 ( .A(n13021), .B(n13022), .Z(n12928) );
  NAND U12825 ( .A(n12730), .B(n12581), .Z(n13020) );
  XOR U12826 ( .A(n12938), .B(n13023), .Z(n12931) );
  IV U12827 ( .A(n12937), .Z(n13023) );
  XNOR U12828 ( .A(n12934), .B(n13024), .Z(n12937) );
  XOR U12829 ( .A(n13025), .B(n13026), .Z(n12934) );
  NANDN U12830 ( .B(n13027), .A(n13028), .Z(n13025) );
  XOR U12831 ( .A(n13026), .B(n13029), .Z(n13028) );
  XOR U12832 ( .A(n12944), .B(n13030), .Z(n12938) );
  IV U12833 ( .A(n12943), .Z(n13030) );
  XNOR U12834 ( .A(n12940), .B(n13031), .Z(n12943) );
  XOR U12835 ( .A(n13032), .B(n13033), .Z(n12940) );
  ANDN U12836 ( .A(n13034), .B(n13035), .Z(n13033) );
  XNOR U12837 ( .A(n13032), .B(n13036), .Z(n13034) );
  XOR U12838 ( .A(n12950), .B(n13037), .Z(n12944) );
  IV U12839 ( .A(n12949), .Z(n13037) );
  XNOR U12840 ( .A(n12946), .B(n13024), .Z(n12949) );
  AND U12841 ( .A(n13181), .B(n12827), .Z(n13024) );
  XOR U12842 ( .A(n13038), .B(n13039), .Z(n12946) );
  ANDN U12843 ( .A(n13040), .B(n13041), .Z(n13039) );
  XNOR U12844 ( .A(n13038), .B(n13042), .Z(n13040) );
  XNOR U12845 ( .A(n12961), .B(n12923), .Z(n12950) );
  NANDN U12846 ( .B(n12845), .A(n12321), .Z(n12923) );
  XNOR U12847 ( .A(n13043), .B(e_input[6]), .Z(n12321) );
  NANDN U12848 ( .B(n12847), .A(n13044), .Z(n13043) );
  XOR U12849 ( .A(n13045), .B(n12956), .Z(n13044) );
  XNOR U12850 ( .A(n12954), .B(n13045), .Z(n12956) );
  XOR U12851 ( .A(n13046), .B(n13047), .Z(n12954) );
  ANDN U12852 ( .A(n13046), .B(n13048), .Z(n13047) );
  IV U12853 ( .A(e_input[6]), .Z(n13045) );
  XNOR U12854 ( .A(n12958), .B(n13049), .Z(n12961) );
  AND U12855 ( .A(n12730), .B(n12581), .Z(n13049) );
  XOR U12856 ( .A(n13050), .B(n13051), .Z(n12958) );
  ANDN U12857 ( .A(n13052), .B(n13053), .Z(n13051) );
  XNOR U12858 ( .A(n13021), .B(n13050), .Z(n13052) );
  XOR U12859 ( .A(n13054), .B(n13013), .Z(n13016) );
  XOR U12860 ( .A(n13055), .B(n13056), .Z(n13013) );
  XNOR U12861 ( .A(n13011), .B(n13014), .Z(n13054) );
  XOR U12862 ( .A(n13057), .B(n12969), .Z(n13011) );
  XOR U12863 ( .A(n12976), .B(n13058), .Z(n12969) );
  IV U12864 ( .A(n12974), .Z(n13058) );
  XNOR U12865 ( .A(n13059), .B(n12973), .Z(n12974) );
  OR U12866 ( .A(n13060), .B(n13061), .Z(n12973) );
  NANDN U12867 ( .B(n6541), .A(n12644), .Z(n13059) );
  XOR U12868 ( .A(n12983), .B(n13062), .Z(n12976) );
  IV U12869 ( .A(n12982), .Z(n13062) );
  XNOR U12870 ( .A(n12979), .B(n13063), .Z(n12982) );
  XOR U12871 ( .A(n13064), .B(n13065), .Z(n12979) );
  NANDN U12872 ( .B(n13066), .A(n13067), .Z(n13064) );
  XOR U12873 ( .A(n13065), .B(n13068), .Z(n13067) );
  XOR U12874 ( .A(n12989), .B(n13069), .Z(n12983) );
  IV U12875 ( .A(n12988), .Z(n13069) );
  XNOR U12876 ( .A(n12985), .B(n13070), .Z(n12988) );
  XOR U12877 ( .A(n13071), .B(n13072), .Z(n12985) );
  ANDN U12878 ( .A(n13073), .B(n13074), .Z(n13072) );
  XNOR U12879 ( .A(n13071), .B(n13075), .Z(n13073) );
  XOR U12880 ( .A(n12995), .B(n13076), .Z(n12989) );
  IV U12881 ( .A(n12994), .Z(n13076) );
  XNOR U12882 ( .A(n12991), .B(n13063), .Z(n12994) );
  AND U12883 ( .A(n13207), .B(n12880), .Z(n13063) );
  XOR U12884 ( .A(n13077), .B(n13078), .Z(n12991) );
  ANDN U12885 ( .A(n13079), .B(n13080), .Z(n13078) );
  XNOR U12886 ( .A(n13077), .B(n13081), .Z(n13079) );
  XNOR U12887 ( .A(n13000), .B(n12968), .Z(n12995) );
  XNOR U12888 ( .A(n12997), .B(n13082), .Z(n13000) );
  AND U12889 ( .A(n6527), .B(n12644), .Z(n13082) );
  XOR U12890 ( .A(n13083), .B(n13084), .Z(n12997) );
  ANDN U12891 ( .A(n13085), .B(n13086), .Z(n13084) );
  XNOR U12892 ( .A(n13060), .B(n13083), .Z(n13085) );
  XOR U12893 ( .A(n13087), .B(n12968), .Z(n13057) );
  NANDN U12894 ( .B(n6808), .A(n12387), .Z(n12968) );
  XOR U12895 ( .A(n13088), .B(n13089), .Z(n12387) );
  AND U12896 ( .A(n6809), .B(n13090), .Z(n13089) );
  XNOR U12897 ( .A(n13088), .B(n13007), .Z(n13090) );
  XOR U12898 ( .A(n13005), .B(n13088), .Z(n13007) );
  XOR U12899 ( .A(n13091), .B(n13092), .Z(n13005) );
  ANDN U12900 ( .A(n13091), .B(n13093), .Z(n13092) );
  XNOR U12901 ( .A(n13094), .B(e_input[23]), .Z(n13088) );
  IV U12902 ( .A(n13009), .Z(n13087) );
  XOR U12903 ( .A(n13095), .B(n13096), .Z(n13009) );
  AND U12904 ( .A(n13097), .B(n13098), .Z(n13096) );
  XNOR U12905 ( .A(n13095), .B(n13099), .Z(n13098) );
  XOR U12906 ( .A(n13100), .B(n13101), .Z(n13014) );
  AND U12907 ( .A(n13102), .B(n13103), .Z(n13101) );
  XNOR U12908 ( .A(n13022), .B(n13104), .Z(n13103) );
  XNOR U12909 ( .A(n13021), .B(n13100), .Z(n13104) );
  XOR U12910 ( .A(n13029), .B(n13105), .Z(n13022) );
  IV U12911 ( .A(n13027), .Z(n13105) );
  XNOR U12912 ( .A(n13106), .B(n13026), .Z(n13027) );
  OR U12913 ( .A(n13107), .B(n13108), .Z(n13026) );
  NAND U12914 ( .A(n12730), .B(n12827), .Z(n13106) );
  XOR U12915 ( .A(n13036), .B(n13109), .Z(n13029) );
  IV U12916 ( .A(n13035), .Z(n13109) );
  XNOR U12917 ( .A(n13032), .B(n13110), .Z(n13035) );
  XOR U12918 ( .A(n13111), .B(n13112), .Z(n13032) );
  NANDN U12919 ( .B(n13113), .A(n13114), .Z(n13111) );
  XOR U12920 ( .A(n13112), .B(n13115), .Z(n13114) );
  XOR U12921 ( .A(n13042), .B(n13116), .Z(n13036) );
  IV U12922 ( .A(n13041), .Z(n13116) );
  XNOR U12923 ( .A(n13038), .B(n13110), .Z(n13041) );
  AND U12924 ( .A(n13181), .B(n13031), .Z(n13110) );
  XNOR U12925 ( .A(n13117), .B(n13118), .Z(n13038) );
  ANDN U12926 ( .A(n13119), .B(n13120), .Z(n13118) );
  XOR U12927 ( .A(n13117), .B(n13121), .Z(n13119) );
  XNOR U12928 ( .A(n13053), .B(n13021), .Z(n13042) );
  NANDN U12929 ( .B(n12845), .A(n12581), .Z(n13021) );
  XNOR U12930 ( .A(n13122), .B(e_input[5]), .Z(n12581) );
  NANDN U12931 ( .B(n12847), .A(n13123), .Z(n13122) );
  XOR U12932 ( .A(n13124), .B(n13048), .Z(n13123) );
  XNOR U12933 ( .A(n13046), .B(n13124), .Z(n13048) );
  XOR U12934 ( .A(n13125), .B(n13126), .Z(n13046) );
  ANDN U12935 ( .A(n13125), .B(n13127), .Z(n13126) );
  IV U12936 ( .A(e_input[5]), .Z(n13124) );
  XNOR U12937 ( .A(n13050), .B(n13128), .Z(n13053) );
  AND U12938 ( .A(n12730), .B(n12827), .Z(n13128) );
  ANDN U12939 ( .A(n13129), .B(n13130), .Z(n13050) );
  NANDN U12940 ( .B(n13131), .A(n13132), .Z(n13129) );
  XOR U12941 ( .A(n13107), .B(n13130), .Z(n13132) );
  XOR U12942 ( .A(n13133), .B(n13099), .Z(n13102) );
  XOR U12943 ( .A(n13134), .B(n13135), .Z(n13099) );
  XNOR U12944 ( .A(n13097), .B(n13100), .Z(n13133) );
  XOR U12945 ( .A(n13136), .B(n13061), .Z(n13097) );
  XOR U12946 ( .A(n13068), .B(n13137), .Z(n13061) );
  IV U12947 ( .A(n13066), .Z(n13137) );
  XNOR U12948 ( .A(n13138), .B(n13065), .Z(n13066) );
  OR U12949 ( .A(n13139), .B(n13140), .Z(n13065) );
  NANDN U12950 ( .B(n6541), .A(n12880), .Z(n13138) );
  XOR U12951 ( .A(n13075), .B(n13141), .Z(n13068) );
  IV U12952 ( .A(n13074), .Z(n13141) );
  XNOR U12953 ( .A(n13071), .B(n13142), .Z(n13074) );
  XOR U12954 ( .A(n13143), .B(n13144), .Z(n13071) );
  NANDN U12955 ( .B(n13145), .A(n13146), .Z(n13143) );
  XOR U12956 ( .A(n13144), .B(n13147), .Z(n13146) );
  XOR U12957 ( .A(n13081), .B(n13148), .Z(n13075) );
  IV U12958 ( .A(n13080), .Z(n13148) );
  XNOR U12959 ( .A(n13077), .B(n13142), .Z(n13080) );
  AND U12960 ( .A(n13207), .B(n13070), .Z(n13142) );
  XOR U12961 ( .A(n13149), .B(n13150), .Z(n13077) );
  ANDN U12962 ( .A(n13151), .B(n13152), .Z(n13150) );
  XNOR U12963 ( .A(n13149), .B(n13153), .Z(n13151) );
  XNOR U12964 ( .A(n13086), .B(n13060), .Z(n13081) );
  XNOR U12965 ( .A(n13083), .B(n13154), .Z(n13086) );
  AND U12966 ( .A(n6527), .B(n12880), .Z(n13154) );
  XOR U12967 ( .A(n13155), .B(n13156), .Z(n13083) );
  ANDN U12968 ( .A(n13157), .B(n13158), .Z(n13156) );
  XNOR U12969 ( .A(n13139), .B(n13155), .Z(n13157) );
  XOR U12970 ( .A(n13159), .B(n13060), .Z(n13136) );
  NANDN U12971 ( .B(n6808), .A(n12644), .Z(n13060) );
  XOR U12972 ( .A(n13160), .B(n13161), .Z(n12644) );
  AND U12973 ( .A(n6809), .B(n13162), .Z(n13161) );
  XNOR U12974 ( .A(n13160), .B(n13093), .Z(n13162) );
  XOR U12975 ( .A(n13091), .B(n13160), .Z(n13093) );
  XOR U12976 ( .A(n13163), .B(n13164), .Z(n13091) );
  ANDN U12977 ( .A(n13163), .B(n13165), .Z(n13164) );
  XNOR U12978 ( .A(n13166), .B(e_input[22]), .Z(n13160) );
  IV U12979 ( .A(n13095), .Z(n13159) );
  XOR U12980 ( .A(n13167), .B(n13168), .Z(n13095) );
  AND U12981 ( .A(n13169), .B(n13170), .Z(n13168) );
  XNOR U12982 ( .A(n13167), .B(n13171), .Z(n13170) );
  XOR U12983 ( .A(n13172), .B(n13173), .Z(n13100) );
  AND U12984 ( .A(n13174), .B(n13175), .Z(n13173) );
  XNOR U12985 ( .A(n13108), .B(n13176), .Z(n13175) );
  XNOR U12986 ( .A(n13107), .B(n13172), .Z(n13176) );
  XOR U12987 ( .A(n13115), .B(n13177), .Z(n13108) );
  IV U12988 ( .A(n13113), .Z(n13177) );
  XNOR U12989 ( .A(n13178), .B(n13112), .Z(n13113) );
  OR U12990 ( .A(n13179), .B(n13180), .Z(n13112) );
  NAND U12991 ( .A(n12730), .B(n13031), .Z(n13178) );
  XNOR U12992 ( .A(n13121), .B(n13120), .Z(n13115) );
  NAND U12993 ( .A(n13181), .B(n13117), .Z(n13120) );
  XNOR U12994 ( .A(n13182), .B(n13183), .Z(n13117) );
  NANDN U12995 ( .B(n13184), .A(n13185), .Z(n13182) );
  XOR U12996 ( .A(n13183), .B(n13186), .Z(n13185) );
  XNOR U12997 ( .A(n13131), .B(n13107), .Z(n13121) );
  NANDN U12998 ( .B(n12845), .A(n12827), .Z(n13107) );
  XNOR U12999 ( .A(n13187), .B(e_input[4]), .Z(n12827) );
  NANDN U13000 ( .B(n12847), .A(n13188), .Z(n13187) );
  XOR U13001 ( .A(n13189), .B(n13127), .Z(n13188) );
  XNOR U13002 ( .A(n13125), .B(n13189), .Z(n13127) );
  XOR U13003 ( .A(n13190), .B(n13191), .Z(n13125) );
  ANDN U13004 ( .A(n13190), .B(n13192), .Z(n13191) );
  IV U13005 ( .A(e_input[4]), .Z(n13189) );
  XOR U13006 ( .A(n13130), .B(n13193), .Z(n13131) );
  AND U13007 ( .A(n12730), .B(n13031), .Z(n13193) );
  NANDN U13008 ( .B(n13194), .A(n13195), .Z(n13130) );
  NANDN U13009 ( .B(n13196), .A(n13197), .Z(n13195) );
  XOR U13010 ( .A(n13194), .B(n13179), .Z(n13197) );
  XOR U13011 ( .A(n13198), .B(n13171), .Z(n13174) );
  XOR U13012 ( .A(n13199), .B(n13200), .Z(n13171) );
  XNOR U13013 ( .A(n13169), .B(n13172), .Z(n13198) );
  XOR U13014 ( .A(n13201), .B(n13140), .Z(n13169) );
  XOR U13015 ( .A(n13147), .B(n13202), .Z(n13140) );
  IV U13016 ( .A(n13145), .Z(n13202) );
  XNOR U13017 ( .A(n13203), .B(n13144), .Z(n13145) );
  OR U13018 ( .A(n13204), .B(n13205), .Z(n13144) );
  NANDN U13019 ( .B(n6541), .A(n13070), .Z(n13203) );
  XOR U13020 ( .A(n13153), .B(n13206), .Z(n13147) );
  IV U13021 ( .A(n13152), .Z(n13206) );
  XNOR U13022 ( .A(n13149), .B(n13207), .Z(n13152) );
  XNOR U13023 ( .A(n13208), .B(n13209), .Z(n13149) );
  NANDN U13024 ( .B(n13210), .A(n13211), .Z(n13208) );
  XNOR U13025 ( .A(n13209), .B(n13212), .Z(n13211) );
  XNOR U13026 ( .A(n13158), .B(n13139), .Z(n13153) );
  XNOR U13027 ( .A(n13155), .B(n13213), .Z(n13158) );
  AND U13028 ( .A(n6527), .B(n13070), .Z(n13213) );
  XOR U13029 ( .A(n13214), .B(n13215), .Z(n13155) );
  ANDN U13030 ( .A(n13216), .B(n13217), .Z(n13215) );
  XNOR U13031 ( .A(n13204), .B(n13214), .Z(n13216) );
  XOR U13032 ( .A(n13218), .B(n13139), .Z(n13201) );
  NANDN U13033 ( .B(n6808), .A(n12880), .Z(n13139) );
  XOR U13034 ( .A(n13219), .B(n13220), .Z(n12880) );
  AND U13035 ( .A(n6809), .B(n13221), .Z(n13220) );
  XNOR U13036 ( .A(n13219), .B(n13165), .Z(n13221) );
  XOR U13037 ( .A(n13163), .B(n13219), .Z(n13165) );
  XOR U13038 ( .A(n13222), .B(n13223), .Z(n13163) );
  ANDN U13039 ( .A(n13222), .B(n13224), .Z(n13223) );
  XNOR U13040 ( .A(n13225), .B(e_input[21]), .Z(n13219) );
  IV U13041 ( .A(n13167), .Z(n13218) );
  XOR U13042 ( .A(n13226), .B(n13227), .Z(n13167) );
  AND U13043 ( .A(n13228), .B(n13229), .Z(n13227) );
  XNOR U13044 ( .A(n13226), .B(n13230), .Z(n13229) );
  XOR U13045 ( .A(n13231), .B(n13232), .Z(n13172) );
  AND U13046 ( .A(n13233), .B(n13234), .Z(n13232) );
  XNOR U13047 ( .A(n13180), .B(n13235), .Z(n13234) );
  XNOR U13048 ( .A(n13179), .B(n13231), .Z(n13235) );
  XOR U13049 ( .A(n13186), .B(n13236), .Z(n13180) );
  IV U13050 ( .A(n13184), .Z(n13236) );
  XNOR U13051 ( .A(n13237), .B(n13183), .Z(n13184) );
  OR U13052 ( .A(n13238), .B(n13239), .Z(n13183) );
  XNOR U13053 ( .A(n13196), .B(n13179), .Z(n13186) );
  NANDN U13054 ( .B(n12845), .A(n13031), .Z(n13179) );
  XNOR U13055 ( .A(n13240), .B(e_input[3]), .Z(n13031) );
  NANDN U13056 ( .B(n12847), .A(n13241), .Z(n13240) );
  XOR U13057 ( .A(n13242), .B(n13192), .Z(n13241) );
  XNOR U13058 ( .A(n13190), .B(n13242), .Z(n13192) );
  XNOR U13059 ( .A(n13243), .B(n13244), .Z(n13190) );
  NOR U13060 ( .A(n13243), .B(n13245), .Z(n13244) );
  IV U13061 ( .A(e_input[3]), .Z(n13242) );
  XNOR U13062 ( .A(n13237), .B(n13194), .Z(n13196) );
  NAND U13063 ( .A(n12730), .B(n13181), .Z(n13237) );
  XOR U13064 ( .A(n13246), .B(n13230), .Z(n13233) );
  XOR U13065 ( .A(n13247), .B(n13248), .Z(n13230) );
  XNOR U13066 ( .A(n13228), .B(n13231), .Z(n13246) );
  XOR U13067 ( .A(n13249), .B(n13205), .Z(n13228) );
  XOR U13068 ( .A(n13212), .B(n13250), .Z(n13205) );
  IV U13069 ( .A(n13210), .Z(n13250) );
  XOR U13070 ( .A(n13251), .B(n13209), .Z(n13210) );
  NOR U13071 ( .A(n13252), .B(n13253), .Z(n13209) );
  NANDN U13072 ( .B(n6541), .A(n13207), .Z(n13251) );
  XNOR U13073 ( .A(n13217), .B(n13204), .Z(n13212) );
  XNOR U13074 ( .A(n13214), .B(n13254), .Z(n13217) );
  AND U13075 ( .A(n6527), .B(n13207), .Z(n13254) );
  XNOR U13076 ( .A(n13255), .B(n13256), .Z(n13214) );
  NANDN U13077 ( .B(n13257), .A(n13258), .Z(n13255) );
  XNOR U13078 ( .A(n13253), .B(n13256), .Z(n13258) );
  XOR U13079 ( .A(n13259), .B(n13204), .Z(n13249) );
  NANDN U13080 ( .B(n6808), .A(n13070), .Z(n13204) );
  XOR U13081 ( .A(n13260), .B(n13261), .Z(n13070) );
  AND U13082 ( .A(n6809), .B(n13262), .Z(n13261) );
  XNOR U13083 ( .A(n13260), .B(n13224), .Z(n13262) );
  XOR U13084 ( .A(n13222), .B(n13260), .Z(n13224) );
  XNOR U13085 ( .A(n13263), .B(n13264), .Z(n13222) );
  NOR U13086 ( .A(n13263), .B(n13265), .Z(n13264) );
  XNOR U13087 ( .A(n13266), .B(e_input[20]), .Z(n13260) );
  IV U13088 ( .A(n13226), .Z(n13259) );
  XOR U13089 ( .A(n13267), .B(n13268), .Z(n13226) );
  AND U13090 ( .A(n13269), .B(n13270), .Z(n13268) );
  XNOR U13091 ( .A(n13267), .B(n13271), .Z(n13270) );
  XNOR U13092 ( .A(n13272), .B(n13273), .Z(n13231) );
  AND U13093 ( .A(n13274), .B(n13275), .Z(n13273) );
  XNOR U13094 ( .A(n13239), .B(n13276), .Z(n13275) );
  XOR U13095 ( .A(n13238), .B(n13272), .Z(n13276) );
  NANDN U13096 ( .B(n12845), .A(n13181), .Z(n13238) );
  XOR U13097 ( .A(n13277), .B(n13278), .Z(n13239) );
  ANDN U13098 ( .A(n13181), .B(n12845), .Z(n13278) );
  XNOR U13099 ( .A(n13279), .B(e_input[2]), .Z(n13181) );
  NANDN U13100 ( .B(n12847), .A(n13280), .Z(n13279) );
  XOR U13101 ( .A(n13281), .B(n13245), .Z(n13280) );
  XOR U13102 ( .A(n13243), .B(n13281), .Z(n13245) );
  XNOR U13103 ( .A(n13282), .B(\MULT3/B__[0] ), .Z(n13243) );
  OR U13104 ( .A(n13283), .B(\MULT3/B__[0] ), .Z(n13282) );
  IV U13105 ( .A(e_input[2]), .Z(n13281) );
  NAND U13106 ( .A(n13284), .B(n12730), .Z(n13277) );
  AND U13107 ( .A(n12730), .B(n13194), .Z(n13284) );
  XOR U13108 ( .A(n13285), .B(n13271), .Z(n13274) );
  XNOR U13109 ( .A(n13286), .B(n13287), .Z(n13271) );
  IV U13110 ( .A(n13288), .Z(n13286) );
  XOR U13111 ( .A(n13269), .B(n13272), .Z(n13285) );
  XNOR U13112 ( .A(n13289), .B(n13290), .Z(n13269) );
  IV U13113 ( .A(n13252), .Z(n13290) );
  XOR U13114 ( .A(n13291), .B(n13253), .Z(n13252) );
  IV U13115 ( .A(n13257), .Z(n13291) );
  XOR U13116 ( .A(n13292), .B(n13256), .Z(n13257) );
  ANDN U13117 ( .A(n13293), .B(n13294), .Z(n13256) );
  NANDN U13118 ( .B(n6541), .A(n6527), .Z(n13292) );
  XNOR U13119 ( .A(n13267), .B(n13253), .Z(n13289) );
  NANDN U13120 ( .B(n6808), .A(n13207), .Z(n13253) );
  XOR U13121 ( .A(n13295), .B(n13296), .Z(n13207) );
  AND U13122 ( .A(n6809), .B(n13297), .Z(n13296) );
  XNOR U13123 ( .A(n13295), .B(n13265), .Z(n13297) );
  XNOR U13124 ( .A(n13263), .B(n13295), .Z(n13265) );
  XNOR U13125 ( .A(n6808), .B(n13298), .Z(n13263) );
  NOR U13126 ( .A(n13299), .B(n13300), .Z(n13298) );
  XNOR U13127 ( .A(n13301), .B(e_input[19]), .Z(n13295) );
  XOR U13128 ( .A(n13302), .B(n13303), .Z(n13267) );
  NANDN U13129 ( .B(n13304), .A(n13305), .Z(n13302) );
  XOR U13130 ( .A(n13303), .B(n13306), .Z(n13305) );
  XNOR U13131 ( .A(n13307), .B(n13308), .Z(n13272) );
  NAND U13132 ( .A(n13309), .B(n13310), .Z(n13307) );
  XNOR U13133 ( .A(n13194), .B(n13311), .Z(n13310) );
  XNOR U13134 ( .A(n13312), .B(n13194), .Z(n13311) );
  NANDN U13135 ( .B(n12845), .A(n12730), .Z(n13194) );
  XNOR U13136 ( .A(n13313), .B(e_input[1]), .Z(n12730) );
  NANDN U13137 ( .B(n12847), .A(n13314), .Z(n13313) );
  XOR U13138 ( .A(n13315), .B(n13283), .Z(n13314) );
  XNOR U13139 ( .A(\MULT3/B__[0] ), .B(e_input[1]), .Z(n13283) );
  IV U13140 ( .A(e_input[1]), .Z(n13315) );
  IV U13141 ( .A(e_input[8]), .Z(n12847) );
  XNOR U13142 ( .A(n13316), .B(n13304), .Z(n13309) );
  XNOR U13143 ( .A(n13317), .B(n13294), .Z(n13304) );
  NANDN U13144 ( .B(n6808), .A(n6527), .Z(n13294) );
  XNOR U13145 ( .A(n13318), .B(n13319), .Z(n6527) );
  IV U13146 ( .A(n13299), .Z(n6808) );
  XNOR U13147 ( .A(n13293), .B(n13303), .Z(n13317) );
  ANDN U13148 ( .A(n13299), .B(n13320), .Z(n13303) );
  AND U13149 ( .A(n13299), .B(n6527), .Z(n13293) );
  XOR U13150 ( .A(n13318), .B(n13319), .Z(n6541) );
  AND U13151 ( .A(n6809), .B(n13321), .Z(n13319) );
  XOR U13152 ( .A(n13318), .B(n13300), .Z(n13321) );
  XNOR U13153 ( .A(n13322), .B(n13299), .Z(n13300) );
  XNOR U13154 ( .A(n13323), .B(n13324), .Z(n6809) );
  AND U13155 ( .A(n13325), .B(n13326), .Z(n13324) );
  XOR U13156 ( .A(n7368), .B(g_input[72]), .Z(n13326) );
  XNOR U13157 ( .A(n7091), .B(n13323), .Z(n13325) );
  XOR U13158 ( .A(n13327), .B(e_input[24]), .Z(n7091) );
  XOR U13159 ( .A(n13328), .B(n13329), .Z(n13323) );
  ANDN U13160 ( .A(n13330), .B(n13327), .Z(n13329) );
  XOR U13161 ( .A(n13328), .B(g_input[72]), .Z(n13327) );
  XNOR U13162 ( .A(n7368), .B(n13328), .Z(n13330) );
  XOR U13163 ( .A(n13331), .B(n13332), .Z(n13328) );
  AND U13164 ( .A(n7367), .B(n13333), .Z(n13332) );
  XNOR U13165 ( .A(n7368), .B(n13331), .Z(n13333) );
  XNOR U13166 ( .A(n13331), .B(g_input[71]), .Z(n7367) );
  XOR U13167 ( .A(n13334), .B(n13335), .Z(n13331) );
  AND U13168 ( .A(n7632), .B(n13336), .Z(n13335) );
  XNOR U13169 ( .A(n7368), .B(n13334), .Z(n13336) );
  XNOR U13170 ( .A(n13334), .B(g_input[70]), .Z(n7632) );
  XOR U13171 ( .A(n13337), .B(n13338), .Z(n13334) );
  AND U13172 ( .A(n7890), .B(n13339), .Z(n13338) );
  XNOR U13173 ( .A(n7368), .B(n13337), .Z(n13339) );
  XNOR U13174 ( .A(n13337), .B(g_input[69]), .Z(n7890) );
  XOR U13175 ( .A(n13340), .B(n13341), .Z(n13337) );
  AND U13176 ( .A(n8141), .B(n13342), .Z(n13341) );
  XNOR U13177 ( .A(n7368), .B(n13340), .Z(n13342) );
  XNOR U13178 ( .A(n13340), .B(g_input[68]), .Z(n8141) );
  XOR U13179 ( .A(n13343), .B(n13344), .Z(n13340) );
  AND U13180 ( .A(n8386), .B(n13345), .Z(n13344) );
  XNOR U13181 ( .A(n7368), .B(n13343), .Z(n13345) );
  XNOR U13182 ( .A(n13343), .B(g_input[67]), .Z(n8386) );
  XOR U13183 ( .A(n13346), .B(n13347), .Z(n13343) );
  AND U13184 ( .A(n8624), .B(n13348), .Z(n13347) );
  XNOR U13185 ( .A(n7368), .B(n13346), .Z(n13348) );
  XNOR U13186 ( .A(n13346), .B(g_input[66]), .Z(n8624) );
  XOR U13187 ( .A(n13349), .B(n13350), .Z(n13346) );
  AND U13188 ( .A(n8856), .B(n13351), .Z(n13350) );
  XNOR U13189 ( .A(n7368), .B(n13349), .Z(n13351) );
  XNOR U13190 ( .A(n13349), .B(g_input[65]), .Z(n8856) );
  XOR U13191 ( .A(n13352), .B(n13353), .Z(n13349) );
  AND U13192 ( .A(n9081), .B(n13354), .Z(n13353) );
  XNOR U13193 ( .A(n7368), .B(n13352), .Z(n13354) );
  XNOR U13194 ( .A(n13352), .B(g_input[64]), .Z(n9081) );
  XOR U13195 ( .A(n13355), .B(n13356), .Z(n13352) );
  AND U13196 ( .A(n9300), .B(n13357), .Z(n13356) );
  XNOR U13197 ( .A(n7368), .B(n13355), .Z(n13357) );
  XNOR U13198 ( .A(n13355), .B(g_input[63]), .Z(n9300) );
  XOR U13199 ( .A(n13358), .B(n13359), .Z(n13355) );
  AND U13200 ( .A(n9512), .B(n13360), .Z(n13359) );
  XNOR U13201 ( .A(n7368), .B(n13358), .Z(n13360) );
  XNOR U13202 ( .A(n13358), .B(g_input[62]), .Z(n9512) );
  XOR U13203 ( .A(n13361), .B(n13362), .Z(n13358) );
  AND U13204 ( .A(n9717), .B(n13363), .Z(n13362) );
  XNOR U13205 ( .A(n7368), .B(n13361), .Z(n13363) );
  XNOR U13206 ( .A(n13361), .B(g_input[61]), .Z(n9717) );
  XOR U13207 ( .A(n13364), .B(n13365), .Z(n13361) );
  AND U13208 ( .A(n9915), .B(n13366), .Z(n13365) );
  XNOR U13209 ( .A(n7368), .B(n13364), .Z(n13366) );
  XNOR U13210 ( .A(n13364), .B(g_input[60]), .Z(n9915) );
  XOR U13211 ( .A(n13367), .B(n13368), .Z(n13364) );
  AND U13212 ( .A(n10107), .B(n13369), .Z(n13368) );
  XNOR U13213 ( .A(n7368), .B(n13367), .Z(n13369) );
  XNOR U13214 ( .A(n13367), .B(g_input[59]), .Z(n10107) );
  XOR U13215 ( .A(n13370), .B(n13371), .Z(n13367) );
  AND U13216 ( .A(n10292), .B(n13372), .Z(n13371) );
  XNOR U13217 ( .A(n7368), .B(n13370), .Z(n13372) );
  XNOR U13218 ( .A(n13370), .B(g_input[58]), .Z(n10292) );
  XOR U13219 ( .A(n13373), .B(n13374), .Z(n13370) );
  AND U13220 ( .A(n10471), .B(n13375), .Z(n13374) );
  XNOR U13221 ( .A(n7368), .B(n13373), .Z(n13375) );
  XNOR U13222 ( .A(n13373), .B(g_input[57]), .Z(n10471) );
  XOR U13223 ( .A(n13376), .B(n13377), .Z(n13373) );
  AND U13224 ( .A(n10643), .B(n13378), .Z(n13377) );
  XNOR U13225 ( .A(n7368), .B(n13376), .Z(n13378) );
  XNOR U13226 ( .A(n13376), .B(g_input[56]), .Z(n10643) );
  XOR U13227 ( .A(n13379), .B(n13380), .Z(n13376) );
  AND U13228 ( .A(n10809), .B(n13381), .Z(n13380) );
  XNOR U13229 ( .A(n7368), .B(n13379), .Z(n13381) );
  XNOR U13230 ( .A(n13379), .B(g_input[55]), .Z(n10809) );
  XOR U13231 ( .A(n13382), .B(n13383), .Z(n13379) );
  AND U13232 ( .A(n10968), .B(n13384), .Z(n13383) );
  XNOR U13233 ( .A(n7368), .B(n13382), .Z(n13384) );
  XNOR U13234 ( .A(n13382), .B(g_input[54]), .Z(n10968) );
  XOR U13235 ( .A(n13385), .B(n13386), .Z(n13382) );
  AND U13236 ( .A(n11121), .B(n13387), .Z(n13386) );
  XNOR U13237 ( .A(n7368), .B(n13385), .Z(n13387) );
  XNOR U13238 ( .A(n13385), .B(g_input[53]), .Z(n11121) );
  XOR U13239 ( .A(n13388), .B(n13389), .Z(n13385) );
  AND U13240 ( .A(n11267), .B(n13390), .Z(n13389) );
  XNOR U13241 ( .A(n7368), .B(n13388), .Z(n13390) );
  XNOR U13242 ( .A(n13388), .B(g_input[52]), .Z(n11267) );
  XOR U13243 ( .A(n13391), .B(n13392), .Z(n13388) );
  AND U13244 ( .A(n11407), .B(n13393), .Z(n13392) );
  XNOR U13245 ( .A(n7368), .B(n13391), .Z(n13393) );
  XNOR U13246 ( .A(n13391), .B(g_input[51]), .Z(n11407) );
  XOR U13247 ( .A(n13394), .B(n13395), .Z(n13391) );
  AND U13248 ( .A(n11540), .B(n13396), .Z(n13395) );
  XNOR U13249 ( .A(n7368), .B(n13394), .Z(n13396) );
  XNOR U13250 ( .A(n13394), .B(g_input[50]), .Z(n11540) );
  XOR U13251 ( .A(n13397), .B(n13398), .Z(n13394) );
  AND U13252 ( .A(n11667), .B(n13399), .Z(n13398) );
  XNOR U13253 ( .A(n7368), .B(n13397), .Z(n13399) );
  XNOR U13254 ( .A(n13397), .B(g_input[49]), .Z(n11667) );
  XOR U13255 ( .A(n13400), .B(n13401), .Z(n13397) );
  AND U13256 ( .A(n11796), .B(n13402), .Z(n13401) );
  XNOR U13257 ( .A(n7368), .B(n13400), .Z(n13402) );
  XNOR U13258 ( .A(n13400), .B(g_input[48]), .Z(n11796) );
  XOR U13259 ( .A(n13403), .B(n13404), .Z(n13400) );
  AND U13260 ( .A(n11923), .B(n13405), .Z(n13404) );
  XNOR U13261 ( .A(n7368), .B(n13403), .Z(n13405) );
  XNOR U13262 ( .A(n13403), .B(g_input[47]), .Z(n11923) );
  XOR U13263 ( .A(n13406), .B(n13407), .Z(n13403) );
  AND U13264 ( .A(n12049), .B(n13408), .Z(n13407) );
  XNOR U13265 ( .A(n7368), .B(n13406), .Z(n13408) );
  XNOR U13266 ( .A(n13406), .B(g_input[46]), .Z(n12049) );
  XOR U13267 ( .A(n13409), .B(n13410), .Z(n13406) );
  AND U13268 ( .A(n12176), .B(n13411), .Z(n13410) );
  XNOR U13269 ( .A(n7368), .B(n13409), .Z(n13411) );
  XNOR U13270 ( .A(n13409), .B(g_input[45]), .Z(n12176) );
  XOR U13271 ( .A(n13412), .B(n13413), .Z(n13409) );
  AND U13272 ( .A(n12302), .B(n13414), .Z(n13413) );
  XNOR U13273 ( .A(n7368), .B(n13412), .Z(n13414) );
  XNOR U13274 ( .A(n13412), .B(g_input[44]), .Z(n12302) );
  XOR U13275 ( .A(n13415), .B(n13416), .Z(n13412) );
  AND U13276 ( .A(n12429), .B(n13417), .Z(n13416) );
  XNOR U13277 ( .A(n7368), .B(n13415), .Z(n13417) );
  XNOR U13278 ( .A(n13415), .B(g_input[43]), .Z(n12429) );
  XOR U13279 ( .A(n13418), .B(n13419), .Z(n13415) );
  AND U13280 ( .A(n12555), .B(n13420), .Z(n13419) );
  XNOR U13281 ( .A(n7368), .B(n13418), .Z(n13420) );
  XNOR U13282 ( .A(n13418), .B(g_input[42]), .Z(n12555) );
  XOR U13283 ( .A(n13421), .B(n13422), .Z(n13418) );
  AND U13284 ( .A(n12680), .B(n13423), .Z(n13422) );
  XNOR U13285 ( .A(n7368), .B(n13421), .Z(n13423) );
  XNOR U13286 ( .A(n13421), .B(g_input[41]), .Z(n12680) );
  XOR U13287 ( .A(n13424), .B(n13425), .Z(n13421) );
  AND U13288 ( .A(n12797), .B(n13426), .Z(n13425) );
  XNOR U13289 ( .A(n7368), .B(n13424), .Z(n13426) );
  XNOR U13290 ( .A(n13424), .B(g_input[40]), .Z(n12797) );
  XOR U13291 ( .A(n13427), .B(n13428), .Z(n13424) );
  AND U13292 ( .A(n12910), .B(n13429), .Z(n13428) );
  XNOR U13293 ( .A(n7368), .B(n13427), .Z(n13429) );
  XNOR U13294 ( .A(n13427), .B(g_input[39]), .Z(n12910) );
  XOR U13295 ( .A(n13430), .B(n13431), .Z(n13427) );
  AND U13296 ( .A(n13008), .B(n13432), .Z(n13431) );
  XNOR U13297 ( .A(n7368), .B(n13430), .Z(n13432) );
  IV U13298 ( .A(e_input[24]), .Z(n7368) );
  XNOR U13299 ( .A(n13430), .B(g_input[38]), .Z(n13008) );
  XOR U13300 ( .A(n13433), .B(n13434), .Z(n13430) );
  AND U13301 ( .A(n13094), .B(n13435), .Z(n13434) );
  XOR U13302 ( .A(e_input[23]), .B(n13433), .Z(n13435) );
  XNOR U13303 ( .A(n13433), .B(g_input[37]), .Z(n13094) );
  XOR U13304 ( .A(n13436), .B(n13437), .Z(n13433) );
  AND U13305 ( .A(n13166), .B(n13438), .Z(n13437) );
  XOR U13306 ( .A(e_input[22]), .B(n13436), .Z(n13438) );
  XNOR U13307 ( .A(n13436), .B(g_input[36]), .Z(n13166) );
  XOR U13308 ( .A(n13439), .B(n13440), .Z(n13436) );
  AND U13309 ( .A(n13225), .B(n13441), .Z(n13440) );
  XOR U13310 ( .A(e_input[21]), .B(n13439), .Z(n13441) );
  XNOR U13311 ( .A(n13439), .B(g_input[35]), .Z(n13225) );
  XOR U13312 ( .A(n13442), .B(n13443), .Z(n13439) );
  AND U13313 ( .A(n13266), .B(n13444), .Z(n13443) );
  XOR U13314 ( .A(e_input[20]), .B(n13442), .Z(n13444) );
  XNOR U13315 ( .A(n13442), .B(g_input[34]), .Z(n13266) );
  XOR U13316 ( .A(n13445), .B(n13446), .Z(n13442) );
  AND U13317 ( .A(n13301), .B(n13447), .Z(n13446) );
  XOR U13318 ( .A(e_input[19]), .B(n13445), .Z(n13447) );
  XNOR U13319 ( .A(n13445), .B(g_input[33]), .Z(n13301) );
  XNOR U13320 ( .A(n13448), .B(n13449), .Z(n13445) );
  NANDN U13321 ( .B(n13450), .A(n13451), .Z(n13448) );
  XOR U13322 ( .A(e_input[18]), .B(n13449), .Z(n13451) );
  IV U13323 ( .A(n13322), .Z(n13318) );
  XOR U13324 ( .A(n13450), .B(e_input[18]), .Z(n13322) );
  XOR U13325 ( .A(n13449), .B(g_input[32]), .Z(n13450) );
  ANDN U13326 ( .A(e_input[17]), .B(g_input[31]), .Z(n13449) );
  XOR U13327 ( .A(n13306), .B(n13308), .Z(n13316) );
  IV U13328 ( .A(n13312), .Z(n13308) );
  NOR U13329 ( .A(n12845), .B(n13452), .Z(n13312) );
  XNOR U13330 ( .A(n13320), .B(n13299), .Z(n13452) );
  XOR U13331 ( .A(e_input[17]), .B(g_input[31]), .Z(n13299) );
  IV U13332 ( .A(\MULT3/B__[0] ), .Z(n12845) );
  XNOR U13333 ( .A(n13453), .B(n13454), .Z(n13306) );
  XOR U13334 ( .A(n13455), .B(n13456), .Z(n2484) );
  IV U13335 ( .A(n13457), .Z(n13456) );
  XOR U13336 ( .A(n13458), .B(n13459), .Z(n2306) );
  IV U13337 ( .A(n13460), .Z(n13459) );
  XOR U13338 ( .A(n13461), .B(n13462), .Z(n2135) );
  IV U13339 ( .A(n13463), .Z(n13462) );
  XOR U13340 ( .A(n13464), .B(n13465), .Z(n1970) );
  IV U13341 ( .A(n13466), .Z(n13465) );
  IV U13342 ( .A(n9), .Z(n794) );
  XNOR U13343 ( .A(n13467), .B(n13468), .Z(n9) );
  ANDN U13344 ( .A(n13469), .B(n13466), .Z(n13468) );
  XNOR U13345 ( .A(n13467), .B(n13470), .Z(n13466) );
  XNOR U13346 ( .A(n13467), .B(n13464), .Z(n13469) );
  XNOR U13347 ( .A(n13471), .B(n13472), .Z(n13464) );
  ANDN U13348 ( .A(n13473), .B(n13474), .Z(n13472) );
  XNOR U13349 ( .A(n13471), .B(n13475), .Z(n13473) );
  XOR U13350 ( .A(n13476), .B(n13477), .Z(n13467) );
  ANDN U13351 ( .A(n13478), .B(n13463), .Z(n13477) );
  XNOR U13352 ( .A(n13476), .B(n13479), .Z(n13463) );
  XNOR U13353 ( .A(n13476), .B(n13461), .Z(n13478) );
  XOR U13354 ( .A(n13475), .B(n13480), .Z(n13461) );
  IV U13355 ( .A(n13474), .Z(n13480) );
  XNOR U13356 ( .A(n13471), .B(n13479), .Z(n13474) );
  AND U13357 ( .A(n13470), .B(n13496), .Z(n13479) );
  XOR U13358 ( .A(n13481), .B(n13482), .Z(n13471) );
  ANDN U13359 ( .A(n13483), .B(n13484), .Z(n13482) );
  XNOR U13360 ( .A(n13481), .B(n13485), .Z(n13483) );
  XNOR U13361 ( .A(n13486), .B(n13487), .Z(n13475) );
  ANDN U13362 ( .A(n13488), .B(n13489), .Z(n13487) );
  XNOR U13363 ( .A(n13486), .B(n13490), .Z(n13488) );
  XOR U13364 ( .A(n13491), .B(n13492), .Z(n13476) );
  ANDN U13365 ( .A(n13493), .B(n13460), .Z(n13492) );
  XNOR U13366 ( .A(n13491), .B(n13494), .Z(n13460) );
  XNOR U13367 ( .A(n13491), .B(n13458), .Z(n13493) );
  XOR U13368 ( .A(n13485), .B(n13495), .Z(n13458) );
  IV U13369 ( .A(n13484), .Z(n13495) );
  XNOR U13370 ( .A(n13481), .B(n13496), .Z(n13484) );
  XOR U13371 ( .A(n13497), .B(n13498), .Z(n13481) );
  ANDN U13372 ( .A(n13499), .B(n13500), .Z(n13498) );
  XNOR U13373 ( .A(n13497), .B(n13501), .Z(n13499) );
  XOR U13374 ( .A(n13490), .B(n13502), .Z(n13485) );
  IV U13375 ( .A(n13489), .Z(n13502) );
  XNOR U13376 ( .A(n13486), .B(n13494), .Z(n13489) );
  AND U13377 ( .A(n13470), .B(n13553), .Z(n13494) );
  XOR U13378 ( .A(n13503), .B(n13504), .Z(n13486) );
  ANDN U13379 ( .A(n13505), .B(n13506), .Z(n13504) );
  XNOR U13380 ( .A(n13503), .B(n13507), .Z(n13505) );
  XNOR U13381 ( .A(n13508), .B(n13509), .Z(n13490) );
  ANDN U13382 ( .A(n13510), .B(n13511), .Z(n13509) );
  XNOR U13383 ( .A(n13508), .B(n13512), .Z(n13510) );
  XOR U13384 ( .A(n13513), .B(n13514), .Z(n13491) );
  ANDN U13385 ( .A(n13515), .B(n13457), .Z(n13514) );
  XNOR U13386 ( .A(n13513), .B(n13516), .Z(n13457) );
  XNOR U13387 ( .A(n13513), .B(n13455), .Z(n13515) );
  XOR U13388 ( .A(n13501), .B(n13517), .Z(n13455) );
  IV U13389 ( .A(n13500), .Z(n13517) );
  XNOR U13390 ( .A(n13497), .B(n13518), .Z(n13500) );
  XOR U13391 ( .A(n13519), .B(n13520), .Z(n13497) );
  ANDN U13392 ( .A(n13521), .B(n13522), .Z(n13520) );
  XNOR U13393 ( .A(n13519), .B(n13523), .Z(n13521) );
  XOR U13394 ( .A(n13507), .B(n13524), .Z(n13501) );
  IV U13395 ( .A(n13506), .Z(n13524) );
  XNOR U13396 ( .A(n13503), .B(n13518), .Z(n13506) );
  AND U13397 ( .A(n13553), .B(n13496), .Z(n13518) );
  XOR U13398 ( .A(n13525), .B(n13526), .Z(n13503) );
  ANDN U13399 ( .A(n13527), .B(n13528), .Z(n13526) );
  XNOR U13400 ( .A(n13525), .B(n13529), .Z(n13527) );
  XOR U13401 ( .A(n13512), .B(n13530), .Z(n13507) );
  IV U13402 ( .A(n13511), .Z(n13530) );
  XNOR U13403 ( .A(n13508), .B(n13516), .Z(n13511) );
  AND U13404 ( .A(n13470), .B(n13636), .Z(n13516) );
  XOR U13405 ( .A(n13531), .B(n13532), .Z(n13508) );
  ANDN U13406 ( .A(n13533), .B(n13534), .Z(n13532) );
  XNOR U13407 ( .A(n13531), .B(n13535), .Z(n13533) );
  XNOR U13408 ( .A(n13536), .B(n13537), .Z(n13512) );
  ANDN U13409 ( .A(n13538), .B(n13539), .Z(n13537) );
  XNOR U13410 ( .A(n13536), .B(n13540), .Z(n13538) );
  XOR U13411 ( .A(n13541), .B(n13542), .Z(n13513) );
  ANDN U13412 ( .A(n13543), .B(n2868), .Z(n13542) );
  XNOR U13413 ( .A(n13541), .B(n13544), .Z(n2868) );
  XNOR U13414 ( .A(n13541), .B(n2866), .Z(n13543) );
  XOR U13415 ( .A(n13523), .B(n13545), .Z(n2866) );
  IV U13416 ( .A(n13522), .Z(n13545) );
  XNOR U13417 ( .A(n13519), .B(n13546), .Z(n13522) );
  XOR U13418 ( .A(n13547), .B(n13548), .Z(n13519) );
  ANDN U13419 ( .A(n13549), .B(n13550), .Z(n13548) );
  XNOR U13420 ( .A(n13547), .B(n13551), .Z(n13549) );
  XOR U13421 ( .A(n13529), .B(n13552), .Z(n13523) );
  IV U13422 ( .A(n13528), .Z(n13552) );
  XNOR U13423 ( .A(n13525), .B(n13553), .Z(n13528) );
  XOR U13424 ( .A(n13554), .B(n13555), .Z(n13525) );
  ANDN U13425 ( .A(n13556), .B(n13557), .Z(n13555) );
  XNOR U13426 ( .A(n13554), .B(n13558), .Z(n13556) );
  XOR U13427 ( .A(n13535), .B(n13559), .Z(n13529) );
  IV U13428 ( .A(n13534), .Z(n13559) );
  XNOR U13429 ( .A(n13531), .B(n13546), .Z(n13534) );
  AND U13430 ( .A(n13636), .B(n13496), .Z(n13546) );
  XOR U13431 ( .A(n13560), .B(n13561), .Z(n13531) );
  ANDN U13432 ( .A(n13562), .B(n13563), .Z(n13561) );
  XNOR U13433 ( .A(n13560), .B(n13564), .Z(n13562) );
  XOR U13434 ( .A(n13540), .B(n13565), .Z(n13535) );
  IV U13435 ( .A(n13539), .Z(n13565) );
  XNOR U13436 ( .A(n13536), .B(n13544), .Z(n13539) );
  AND U13437 ( .A(n13470), .B(n13745), .Z(n13544) );
  XOR U13438 ( .A(n13566), .B(n13567), .Z(n13536) );
  ANDN U13439 ( .A(n13568), .B(n13569), .Z(n13567) );
  XNOR U13440 ( .A(n13566), .B(n13570), .Z(n13568) );
  XNOR U13441 ( .A(n13571), .B(n13572), .Z(n13540) );
  ANDN U13442 ( .A(n13573), .B(n13574), .Z(n13572) );
  XNOR U13443 ( .A(n13571), .B(n13575), .Z(n13573) );
  XOR U13444 ( .A(n13576), .B(n13577), .Z(n13541) );
  ANDN U13445 ( .A(n13578), .B(n3068), .Z(n13577) );
  XNOR U13446 ( .A(n13576), .B(n13579), .Z(n3068) );
  XNOR U13447 ( .A(n13576), .B(n3066), .Z(n13578) );
  XOR U13448 ( .A(n13551), .B(n13580), .Z(n3066) );
  IV U13449 ( .A(n13550), .Z(n13580) );
  XNOR U13450 ( .A(n13547), .B(n13581), .Z(n13550) );
  XOR U13451 ( .A(n13582), .B(n13583), .Z(n13547) );
  ANDN U13452 ( .A(n13584), .B(n13585), .Z(n13583) );
  XNOR U13453 ( .A(n13582), .B(n13586), .Z(n13584) );
  XOR U13454 ( .A(n13558), .B(n13587), .Z(n13551) );
  IV U13455 ( .A(n13557), .Z(n13587) );
  XNOR U13456 ( .A(n13554), .B(n13588), .Z(n13557) );
  XOR U13457 ( .A(n13589), .B(n13590), .Z(n13554) );
  ANDN U13458 ( .A(n13591), .B(n13592), .Z(n13590) );
  XNOR U13459 ( .A(n13589), .B(n13593), .Z(n13591) );
  XOR U13460 ( .A(n13564), .B(n13594), .Z(n13558) );
  IV U13461 ( .A(n13563), .Z(n13594) );
  XNOR U13462 ( .A(n13560), .B(n13588), .Z(n13563) );
  AND U13463 ( .A(n13636), .B(n13553), .Z(n13588) );
  XOR U13464 ( .A(n13595), .B(n13596), .Z(n13560) );
  ANDN U13465 ( .A(n13597), .B(n13598), .Z(n13596) );
  XNOR U13466 ( .A(n13595), .B(n13599), .Z(n13597) );
  XOR U13467 ( .A(n13570), .B(n13600), .Z(n13564) );
  IV U13468 ( .A(n13569), .Z(n13600) );
  XNOR U13469 ( .A(n13566), .B(n13581), .Z(n13569) );
  AND U13470 ( .A(n13745), .B(n13496), .Z(n13581) );
  XOR U13471 ( .A(n13601), .B(n13602), .Z(n13566) );
  ANDN U13472 ( .A(n13603), .B(n13604), .Z(n13602) );
  XNOR U13473 ( .A(n13601), .B(n13605), .Z(n13603) );
  XOR U13474 ( .A(n13575), .B(n13606), .Z(n13570) );
  IV U13475 ( .A(n13574), .Z(n13606) );
  XNOR U13476 ( .A(n13571), .B(n13579), .Z(n13574) );
  AND U13477 ( .A(n13470), .B(n13880), .Z(n13579) );
  XOR U13478 ( .A(n13607), .B(n13608), .Z(n13571) );
  ANDN U13479 ( .A(n13609), .B(n13610), .Z(n13608) );
  XNOR U13480 ( .A(n13607), .B(n13611), .Z(n13609) );
  XNOR U13481 ( .A(n13612), .B(n13613), .Z(n13575) );
  ANDN U13482 ( .A(n13614), .B(n13615), .Z(n13613) );
  XNOR U13483 ( .A(n13612), .B(n13616), .Z(n13614) );
  XOR U13484 ( .A(n13617), .B(n13618), .Z(n13576) );
  ANDN U13485 ( .A(n13619), .B(n3275), .Z(n13618) );
  XNOR U13486 ( .A(n13617), .B(n13620), .Z(n3275) );
  XNOR U13487 ( .A(n13617), .B(n3273), .Z(n13619) );
  XOR U13488 ( .A(n13586), .B(n13621), .Z(n3273) );
  IV U13489 ( .A(n13585), .Z(n13621) );
  XNOR U13490 ( .A(n13582), .B(n13622), .Z(n13585) );
  XOR U13491 ( .A(n13623), .B(n13624), .Z(n13582) );
  ANDN U13492 ( .A(n13625), .B(n13626), .Z(n13624) );
  XNOR U13493 ( .A(n13623), .B(n13627), .Z(n13625) );
  XOR U13494 ( .A(n13593), .B(n13628), .Z(n13586) );
  IV U13495 ( .A(n13592), .Z(n13628) );
  XNOR U13496 ( .A(n13589), .B(n13629), .Z(n13592) );
  XOR U13497 ( .A(n13630), .B(n13631), .Z(n13589) );
  ANDN U13498 ( .A(n13632), .B(n13633), .Z(n13631) );
  XNOR U13499 ( .A(n13630), .B(n13634), .Z(n13632) );
  XOR U13500 ( .A(n13599), .B(n13635), .Z(n13593) );
  IV U13501 ( .A(n13598), .Z(n13635) );
  XNOR U13502 ( .A(n13595), .B(n13636), .Z(n13598) );
  XOR U13503 ( .A(n13637), .B(n13638), .Z(n13595) );
  ANDN U13504 ( .A(n13639), .B(n13640), .Z(n13638) );
  XNOR U13505 ( .A(n13637), .B(n13641), .Z(n13639) );
  XOR U13506 ( .A(n13605), .B(n13642), .Z(n13599) );
  IV U13507 ( .A(n13604), .Z(n13642) );
  XNOR U13508 ( .A(n13601), .B(n13629), .Z(n13604) );
  AND U13509 ( .A(n13745), .B(n13553), .Z(n13629) );
  XOR U13510 ( .A(n13643), .B(n13644), .Z(n13601) );
  ANDN U13511 ( .A(n13645), .B(n13646), .Z(n13644) );
  XNOR U13512 ( .A(n13643), .B(n13647), .Z(n13645) );
  XOR U13513 ( .A(n13611), .B(n13648), .Z(n13605) );
  IV U13514 ( .A(n13610), .Z(n13648) );
  XNOR U13515 ( .A(n13607), .B(n13622), .Z(n13610) );
  AND U13516 ( .A(n13880), .B(n13496), .Z(n13622) );
  XOR U13517 ( .A(n13649), .B(n13650), .Z(n13607) );
  ANDN U13518 ( .A(n13651), .B(n13652), .Z(n13650) );
  XNOR U13519 ( .A(n13649), .B(n13653), .Z(n13651) );
  XOR U13520 ( .A(n13616), .B(n13654), .Z(n13611) );
  IV U13521 ( .A(n13615), .Z(n13654) );
  XNOR U13522 ( .A(n13612), .B(n13620), .Z(n13615) );
  AND U13523 ( .A(n13470), .B(n14041), .Z(n13620) );
  XOR U13524 ( .A(n13655), .B(n13656), .Z(n13612) );
  ANDN U13525 ( .A(n13657), .B(n13658), .Z(n13656) );
  XNOR U13526 ( .A(n13655), .B(n13659), .Z(n13657) );
  XNOR U13527 ( .A(n13660), .B(n13661), .Z(n13616) );
  ANDN U13528 ( .A(n13662), .B(n13663), .Z(n13661) );
  XNOR U13529 ( .A(n13660), .B(n13664), .Z(n13662) );
  XOR U13530 ( .A(n13665), .B(n13666), .Z(n13617) );
  ANDN U13531 ( .A(n13667), .B(n3488), .Z(n13666) );
  XNOR U13532 ( .A(n13665), .B(n13668), .Z(n3488) );
  XNOR U13533 ( .A(n13665), .B(n3486), .Z(n13667) );
  XOR U13534 ( .A(n13627), .B(n13669), .Z(n3486) );
  IV U13535 ( .A(n13626), .Z(n13669) );
  XNOR U13536 ( .A(n13623), .B(n13670), .Z(n13626) );
  XOR U13537 ( .A(n13671), .B(n13672), .Z(n13623) );
  ANDN U13538 ( .A(n13673), .B(n13674), .Z(n13672) );
  XNOR U13539 ( .A(n13671), .B(n13675), .Z(n13673) );
  XOR U13540 ( .A(n13634), .B(n13676), .Z(n13627) );
  IV U13541 ( .A(n13633), .Z(n13676) );
  XNOR U13542 ( .A(n13630), .B(n13677), .Z(n13633) );
  XOR U13543 ( .A(n13678), .B(n13679), .Z(n13630) );
  ANDN U13544 ( .A(n13680), .B(n13681), .Z(n13679) );
  XNOR U13545 ( .A(n13678), .B(n13682), .Z(n13680) );
  XOR U13546 ( .A(n13641), .B(n13683), .Z(n13634) );
  IV U13547 ( .A(n13640), .Z(n13683) );
  XNOR U13548 ( .A(n13637), .B(n13684), .Z(n13640) );
  XOR U13549 ( .A(n13685), .B(n13686), .Z(n13637) );
  ANDN U13550 ( .A(n13687), .B(n13688), .Z(n13686) );
  XNOR U13551 ( .A(n13685), .B(n13689), .Z(n13687) );
  XOR U13552 ( .A(n13647), .B(n13690), .Z(n13641) );
  IV U13553 ( .A(n13646), .Z(n13690) );
  XNOR U13554 ( .A(n13643), .B(n13684), .Z(n13646) );
  AND U13555 ( .A(n13745), .B(n13636), .Z(n13684) );
  XOR U13556 ( .A(n13691), .B(n13692), .Z(n13643) );
  ANDN U13557 ( .A(n13693), .B(n13694), .Z(n13692) );
  XNOR U13558 ( .A(n13691), .B(n13695), .Z(n13693) );
  XOR U13559 ( .A(n13653), .B(n13696), .Z(n13647) );
  IV U13560 ( .A(n13652), .Z(n13696) );
  XNOR U13561 ( .A(n13649), .B(n13677), .Z(n13652) );
  AND U13562 ( .A(n13880), .B(n13553), .Z(n13677) );
  XOR U13563 ( .A(n13697), .B(n13698), .Z(n13649) );
  ANDN U13564 ( .A(n13699), .B(n13700), .Z(n13698) );
  XNOR U13565 ( .A(n13697), .B(n13701), .Z(n13699) );
  XOR U13566 ( .A(n13659), .B(n13702), .Z(n13653) );
  IV U13567 ( .A(n13658), .Z(n13702) );
  XNOR U13568 ( .A(n13655), .B(n13670), .Z(n13658) );
  AND U13569 ( .A(n14041), .B(n13496), .Z(n13670) );
  XOR U13570 ( .A(n13703), .B(n13704), .Z(n13655) );
  ANDN U13571 ( .A(n13705), .B(n13706), .Z(n13704) );
  XNOR U13572 ( .A(n13703), .B(n13707), .Z(n13705) );
  XOR U13573 ( .A(n13664), .B(n13708), .Z(n13659) );
  IV U13574 ( .A(n13663), .Z(n13708) );
  XNOR U13575 ( .A(n13660), .B(n13668), .Z(n13663) );
  AND U13576 ( .A(n13470), .B(n14228), .Z(n13668) );
  XOR U13577 ( .A(n13709), .B(n13710), .Z(n13660) );
  ANDN U13578 ( .A(n13711), .B(n13712), .Z(n13710) );
  XNOR U13579 ( .A(n13709), .B(n13713), .Z(n13711) );
  XNOR U13580 ( .A(n13714), .B(n13715), .Z(n13664) );
  ANDN U13581 ( .A(n13716), .B(n13717), .Z(n13715) );
  XNOR U13582 ( .A(n13714), .B(n13718), .Z(n13716) );
  XOR U13583 ( .A(n13719), .B(n13720), .Z(n13665) );
  ANDN U13584 ( .A(n13721), .B(n3708), .Z(n13720) );
  XNOR U13585 ( .A(n13719), .B(n13722), .Z(n3708) );
  XNOR U13586 ( .A(n13719), .B(n3706), .Z(n13721) );
  XOR U13587 ( .A(n13675), .B(n13723), .Z(n3706) );
  IV U13588 ( .A(n13674), .Z(n13723) );
  XNOR U13589 ( .A(n13671), .B(n13724), .Z(n13674) );
  XOR U13590 ( .A(n13725), .B(n13726), .Z(n13671) );
  ANDN U13591 ( .A(n13727), .B(n13728), .Z(n13726) );
  XNOR U13592 ( .A(n13725), .B(n13729), .Z(n13727) );
  XOR U13593 ( .A(n13682), .B(n13730), .Z(n13675) );
  IV U13594 ( .A(n13681), .Z(n13730) );
  XNOR U13595 ( .A(n13678), .B(n13731), .Z(n13681) );
  XOR U13596 ( .A(n13732), .B(n13733), .Z(n13678) );
  ANDN U13597 ( .A(n13734), .B(n13735), .Z(n13733) );
  XNOR U13598 ( .A(n13732), .B(n13736), .Z(n13734) );
  XOR U13599 ( .A(n13689), .B(n13737), .Z(n13682) );
  IV U13600 ( .A(n13688), .Z(n13737) );
  XNOR U13601 ( .A(n13685), .B(n13738), .Z(n13688) );
  XOR U13602 ( .A(n13739), .B(n13740), .Z(n13685) );
  ANDN U13603 ( .A(n13741), .B(n13742), .Z(n13740) );
  XNOR U13604 ( .A(n13739), .B(n13743), .Z(n13741) );
  XOR U13605 ( .A(n13695), .B(n13744), .Z(n13689) );
  IV U13606 ( .A(n13694), .Z(n13744) );
  XNOR U13607 ( .A(n13691), .B(n13745), .Z(n13694) );
  XOR U13608 ( .A(n13746), .B(n13747), .Z(n13691) );
  ANDN U13609 ( .A(n13748), .B(n13749), .Z(n13747) );
  XNOR U13610 ( .A(n13746), .B(n13750), .Z(n13748) );
  XOR U13611 ( .A(n13701), .B(n13751), .Z(n13695) );
  IV U13612 ( .A(n13700), .Z(n13751) );
  XNOR U13613 ( .A(n13697), .B(n13738), .Z(n13700) );
  AND U13614 ( .A(n13880), .B(n13636), .Z(n13738) );
  XOR U13615 ( .A(n13752), .B(n13753), .Z(n13697) );
  ANDN U13616 ( .A(n13754), .B(n13755), .Z(n13753) );
  XNOR U13617 ( .A(n13752), .B(n13756), .Z(n13754) );
  XOR U13618 ( .A(n13707), .B(n13757), .Z(n13701) );
  IV U13619 ( .A(n13706), .Z(n13757) );
  XNOR U13620 ( .A(n13703), .B(n13731), .Z(n13706) );
  AND U13621 ( .A(n14041), .B(n13553), .Z(n13731) );
  XOR U13622 ( .A(n13758), .B(n13759), .Z(n13703) );
  ANDN U13623 ( .A(n13760), .B(n13761), .Z(n13759) );
  XNOR U13624 ( .A(n13758), .B(n13762), .Z(n13760) );
  XOR U13625 ( .A(n13713), .B(n13763), .Z(n13707) );
  IV U13626 ( .A(n13712), .Z(n13763) );
  XNOR U13627 ( .A(n13709), .B(n13724), .Z(n13712) );
  AND U13628 ( .A(n14228), .B(n13496), .Z(n13724) );
  XOR U13629 ( .A(n13764), .B(n13765), .Z(n13709) );
  ANDN U13630 ( .A(n13766), .B(n13767), .Z(n13765) );
  XNOR U13631 ( .A(n13764), .B(n13768), .Z(n13766) );
  XOR U13632 ( .A(n13718), .B(n13769), .Z(n13713) );
  IV U13633 ( .A(n13717), .Z(n13769) );
  XNOR U13634 ( .A(n13714), .B(n13722), .Z(n13717) );
  AND U13635 ( .A(n13470), .B(n14441), .Z(n13722) );
  XOR U13636 ( .A(n13770), .B(n13771), .Z(n13714) );
  ANDN U13637 ( .A(n13772), .B(n13773), .Z(n13771) );
  XNOR U13638 ( .A(n13770), .B(n13774), .Z(n13772) );
  XNOR U13639 ( .A(n13775), .B(n13776), .Z(n13718) );
  ANDN U13640 ( .A(n13777), .B(n13778), .Z(n13776) );
  XNOR U13641 ( .A(n13775), .B(n13779), .Z(n13777) );
  XOR U13642 ( .A(n13780), .B(n13781), .Z(n13719) );
  ANDN U13643 ( .A(n13782), .B(n3934), .Z(n13781) );
  XNOR U13644 ( .A(n13780), .B(n13783), .Z(n3934) );
  XNOR U13645 ( .A(n13780), .B(n3932), .Z(n13782) );
  XOR U13646 ( .A(n13729), .B(n13784), .Z(n3932) );
  IV U13647 ( .A(n13728), .Z(n13784) );
  XNOR U13648 ( .A(n13725), .B(n13785), .Z(n13728) );
  XOR U13649 ( .A(n13786), .B(n13787), .Z(n13725) );
  ANDN U13650 ( .A(n13788), .B(n13789), .Z(n13787) );
  XNOR U13651 ( .A(n13786), .B(n13790), .Z(n13788) );
  XOR U13652 ( .A(n13736), .B(n13791), .Z(n13729) );
  IV U13653 ( .A(n13735), .Z(n13791) );
  XNOR U13654 ( .A(n13732), .B(n13792), .Z(n13735) );
  XOR U13655 ( .A(n13793), .B(n13794), .Z(n13732) );
  ANDN U13656 ( .A(n13795), .B(n13796), .Z(n13794) );
  XNOR U13657 ( .A(n13793), .B(n13797), .Z(n13795) );
  XOR U13658 ( .A(n13743), .B(n13798), .Z(n13736) );
  IV U13659 ( .A(n13742), .Z(n13798) );
  XNOR U13660 ( .A(n13739), .B(n13799), .Z(n13742) );
  XOR U13661 ( .A(n13800), .B(n13801), .Z(n13739) );
  ANDN U13662 ( .A(n13802), .B(n13803), .Z(n13801) );
  XNOR U13663 ( .A(n13800), .B(n13804), .Z(n13802) );
  XOR U13664 ( .A(n13750), .B(n13805), .Z(n13743) );
  IV U13665 ( .A(n13749), .Z(n13805) );
  XNOR U13666 ( .A(n13746), .B(n13806), .Z(n13749) );
  XOR U13667 ( .A(n13807), .B(n13808), .Z(n13746) );
  ANDN U13668 ( .A(n13809), .B(n13810), .Z(n13808) );
  XNOR U13669 ( .A(n13807), .B(n13811), .Z(n13809) );
  XOR U13670 ( .A(n13756), .B(n13812), .Z(n13750) );
  IV U13671 ( .A(n13755), .Z(n13812) );
  XNOR U13672 ( .A(n13752), .B(n13806), .Z(n13755) );
  AND U13673 ( .A(n13880), .B(n13745), .Z(n13806) );
  XOR U13674 ( .A(n13813), .B(n13814), .Z(n13752) );
  ANDN U13675 ( .A(n13815), .B(n13816), .Z(n13814) );
  XNOR U13676 ( .A(n13813), .B(n13817), .Z(n13815) );
  XOR U13677 ( .A(n13762), .B(n13818), .Z(n13756) );
  IV U13678 ( .A(n13761), .Z(n13818) );
  XNOR U13679 ( .A(n13758), .B(n13799), .Z(n13761) );
  AND U13680 ( .A(n14041), .B(n13636), .Z(n13799) );
  XOR U13681 ( .A(n13819), .B(n13820), .Z(n13758) );
  ANDN U13682 ( .A(n13821), .B(n13822), .Z(n13820) );
  XNOR U13683 ( .A(n13819), .B(n13823), .Z(n13821) );
  XOR U13684 ( .A(n13768), .B(n13824), .Z(n13762) );
  IV U13685 ( .A(n13767), .Z(n13824) );
  XNOR U13686 ( .A(n13764), .B(n13792), .Z(n13767) );
  AND U13687 ( .A(n14228), .B(n13553), .Z(n13792) );
  XOR U13688 ( .A(n13825), .B(n13826), .Z(n13764) );
  ANDN U13689 ( .A(n13827), .B(n13828), .Z(n13826) );
  XNOR U13690 ( .A(n13825), .B(n13829), .Z(n13827) );
  XOR U13691 ( .A(n13774), .B(n13830), .Z(n13768) );
  IV U13692 ( .A(n13773), .Z(n13830) );
  XNOR U13693 ( .A(n13770), .B(n13785), .Z(n13773) );
  AND U13694 ( .A(n14441), .B(n13496), .Z(n13785) );
  XOR U13695 ( .A(n13831), .B(n13832), .Z(n13770) );
  ANDN U13696 ( .A(n13833), .B(n13834), .Z(n13832) );
  XNOR U13697 ( .A(n13831), .B(n13835), .Z(n13833) );
  XOR U13698 ( .A(n13779), .B(n13836), .Z(n13774) );
  IV U13699 ( .A(n13778), .Z(n13836) );
  XNOR U13700 ( .A(n13775), .B(n13783), .Z(n13778) );
  AND U13701 ( .A(n13470), .B(n14680), .Z(n13783) );
  XOR U13702 ( .A(n13837), .B(n13838), .Z(n13775) );
  ANDN U13703 ( .A(n13839), .B(n13840), .Z(n13838) );
  XNOR U13704 ( .A(n13837), .B(n13841), .Z(n13839) );
  XNOR U13705 ( .A(n13842), .B(n13843), .Z(n13779) );
  ANDN U13706 ( .A(n13844), .B(n13845), .Z(n13843) );
  XNOR U13707 ( .A(n13842), .B(n13846), .Z(n13844) );
  XOR U13708 ( .A(n13847), .B(n13848), .Z(n13780) );
  ANDN U13709 ( .A(n13849), .B(n4167), .Z(n13848) );
  XNOR U13710 ( .A(n13847), .B(n13850), .Z(n4167) );
  XNOR U13711 ( .A(n13847), .B(n4165), .Z(n13849) );
  XOR U13712 ( .A(n13790), .B(n13851), .Z(n4165) );
  IV U13713 ( .A(n13789), .Z(n13851) );
  XNOR U13714 ( .A(n13786), .B(n13852), .Z(n13789) );
  XOR U13715 ( .A(n13853), .B(n13854), .Z(n13786) );
  ANDN U13716 ( .A(n13855), .B(n13856), .Z(n13854) );
  XNOR U13717 ( .A(n13853), .B(n13857), .Z(n13855) );
  XOR U13718 ( .A(n13797), .B(n13858), .Z(n13790) );
  IV U13719 ( .A(n13796), .Z(n13858) );
  XNOR U13720 ( .A(n13793), .B(n13859), .Z(n13796) );
  XOR U13721 ( .A(n13860), .B(n13861), .Z(n13793) );
  ANDN U13722 ( .A(n13862), .B(n13863), .Z(n13861) );
  XNOR U13723 ( .A(n13860), .B(n13864), .Z(n13862) );
  XOR U13724 ( .A(n13804), .B(n13865), .Z(n13797) );
  IV U13725 ( .A(n13803), .Z(n13865) );
  XNOR U13726 ( .A(n13800), .B(n13866), .Z(n13803) );
  XOR U13727 ( .A(n13867), .B(n13868), .Z(n13800) );
  ANDN U13728 ( .A(n13869), .B(n13870), .Z(n13868) );
  XNOR U13729 ( .A(n13867), .B(n13871), .Z(n13869) );
  XOR U13730 ( .A(n13811), .B(n13872), .Z(n13804) );
  IV U13731 ( .A(n13810), .Z(n13872) );
  XNOR U13732 ( .A(n13807), .B(n13873), .Z(n13810) );
  XOR U13733 ( .A(n13874), .B(n13875), .Z(n13807) );
  ANDN U13734 ( .A(n13876), .B(n13877), .Z(n13875) );
  XNOR U13735 ( .A(n13874), .B(n13878), .Z(n13876) );
  XOR U13736 ( .A(n13817), .B(n13879), .Z(n13811) );
  IV U13737 ( .A(n13816), .Z(n13879) );
  XNOR U13738 ( .A(n13813), .B(n13880), .Z(n13816) );
  XOR U13739 ( .A(n13881), .B(n13882), .Z(n13813) );
  ANDN U13740 ( .A(n13883), .B(n13884), .Z(n13882) );
  XNOR U13741 ( .A(n13881), .B(n13885), .Z(n13883) );
  XOR U13742 ( .A(n13823), .B(n13886), .Z(n13817) );
  IV U13743 ( .A(n13822), .Z(n13886) );
  XNOR U13744 ( .A(n13819), .B(n13873), .Z(n13822) );
  AND U13745 ( .A(n14041), .B(n13745), .Z(n13873) );
  XOR U13746 ( .A(n13887), .B(n13888), .Z(n13819) );
  ANDN U13747 ( .A(n13889), .B(n13890), .Z(n13888) );
  XNOR U13748 ( .A(n13887), .B(n13891), .Z(n13889) );
  XOR U13749 ( .A(n13829), .B(n13892), .Z(n13823) );
  IV U13750 ( .A(n13828), .Z(n13892) );
  XNOR U13751 ( .A(n13825), .B(n13866), .Z(n13828) );
  AND U13752 ( .A(n14228), .B(n13636), .Z(n13866) );
  XOR U13753 ( .A(n13893), .B(n13894), .Z(n13825) );
  ANDN U13754 ( .A(n13895), .B(n13896), .Z(n13894) );
  XNOR U13755 ( .A(n13893), .B(n13897), .Z(n13895) );
  XOR U13756 ( .A(n13835), .B(n13898), .Z(n13829) );
  IV U13757 ( .A(n13834), .Z(n13898) );
  XNOR U13758 ( .A(n13831), .B(n13859), .Z(n13834) );
  AND U13759 ( .A(n14441), .B(n13553), .Z(n13859) );
  XOR U13760 ( .A(n13899), .B(n13900), .Z(n13831) );
  ANDN U13761 ( .A(n13901), .B(n13902), .Z(n13900) );
  XNOR U13762 ( .A(n13899), .B(n13903), .Z(n13901) );
  XOR U13763 ( .A(n13841), .B(n13904), .Z(n13835) );
  IV U13764 ( .A(n13840), .Z(n13904) );
  XNOR U13765 ( .A(n13837), .B(n13852), .Z(n13840) );
  AND U13766 ( .A(n14680), .B(n13496), .Z(n13852) );
  XOR U13767 ( .A(n13905), .B(n13906), .Z(n13837) );
  ANDN U13768 ( .A(n13907), .B(n13908), .Z(n13906) );
  XNOR U13769 ( .A(n13905), .B(n13909), .Z(n13907) );
  XOR U13770 ( .A(n13846), .B(n13910), .Z(n13841) );
  IV U13771 ( .A(n13845), .Z(n13910) );
  XNOR U13772 ( .A(n13842), .B(n13850), .Z(n13845) );
  AND U13773 ( .A(n13470), .B(n14945), .Z(n13850) );
  XOR U13774 ( .A(n13911), .B(n13912), .Z(n13842) );
  ANDN U13775 ( .A(n13913), .B(n13914), .Z(n13912) );
  XNOR U13776 ( .A(n13911), .B(n13915), .Z(n13913) );
  XNOR U13777 ( .A(n13916), .B(n13917), .Z(n13846) );
  ANDN U13778 ( .A(n13918), .B(n13919), .Z(n13917) );
  XNOR U13779 ( .A(n13916), .B(n13920), .Z(n13918) );
  XOR U13780 ( .A(n13921), .B(n13922), .Z(n13847) );
  ANDN U13781 ( .A(n13923), .B(n4406), .Z(n13922) );
  XNOR U13782 ( .A(n13921), .B(n13924), .Z(n4406) );
  XNOR U13783 ( .A(n13921), .B(n4404), .Z(n13923) );
  XOR U13784 ( .A(n13857), .B(n13925), .Z(n4404) );
  IV U13785 ( .A(n13856), .Z(n13925) );
  XNOR U13786 ( .A(n13853), .B(n13926), .Z(n13856) );
  XOR U13787 ( .A(n13927), .B(n13928), .Z(n13853) );
  ANDN U13788 ( .A(n13929), .B(n13930), .Z(n13928) );
  XNOR U13789 ( .A(n13927), .B(n13931), .Z(n13929) );
  XOR U13790 ( .A(n13864), .B(n13932), .Z(n13857) );
  IV U13791 ( .A(n13863), .Z(n13932) );
  XNOR U13792 ( .A(n13860), .B(n13933), .Z(n13863) );
  XOR U13793 ( .A(n13934), .B(n13935), .Z(n13860) );
  ANDN U13794 ( .A(n13936), .B(n13937), .Z(n13935) );
  XNOR U13795 ( .A(n13934), .B(n13938), .Z(n13936) );
  XOR U13796 ( .A(n13871), .B(n13939), .Z(n13864) );
  IV U13797 ( .A(n13870), .Z(n13939) );
  XNOR U13798 ( .A(n13867), .B(n13940), .Z(n13870) );
  XOR U13799 ( .A(n13941), .B(n13942), .Z(n13867) );
  ANDN U13800 ( .A(n13943), .B(n13944), .Z(n13942) );
  XNOR U13801 ( .A(n13941), .B(n13945), .Z(n13943) );
  XOR U13802 ( .A(n13878), .B(n13946), .Z(n13871) );
  IV U13803 ( .A(n13877), .Z(n13946) );
  XNOR U13804 ( .A(n13874), .B(n13947), .Z(n13877) );
  XOR U13805 ( .A(n13948), .B(n13949), .Z(n13874) );
  ANDN U13806 ( .A(n13950), .B(n13951), .Z(n13949) );
  XNOR U13807 ( .A(n13948), .B(n13952), .Z(n13950) );
  XOR U13808 ( .A(n13885), .B(n13953), .Z(n13878) );
  IV U13809 ( .A(n13884), .Z(n13953) );
  XNOR U13810 ( .A(n13881), .B(n13954), .Z(n13884) );
  XOR U13811 ( .A(n13955), .B(n13956), .Z(n13881) );
  ANDN U13812 ( .A(n13957), .B(n13958), .Z(n13956) );
  XNOR U13813 ( .A(n13955), .B(n13959), .Z(n13957) );
  XOR U13814 ( .A(n13891), .B(n13960), .Z(n13885) );
  IV U13815 ( .A(n13890), .Z(n13960) );
  XNOR U13816 ( .A(n13887), .B(n13954), .Z(n13890) );
  AND U13817 ( .A(n14041), .B(n13880), .Z(n13954) );
  XOR U13818 ( .A(n13961), .B(n13962), .Z(n13887) );
  ANDN U13819 ( .A(n13963), .B(n13964), .Z(n13962) );
  XNOR U13820 ( .A(n13961), .B(n13965), .Z(n13963) );
  XOR U13821 ( .A(n13897), .B(n13966), .Z(n13891) );
  IV U13822 ( .A(n13896), .Z(n13966) );
  XNOR U13823 ( .A(n13893), .B(n13947), .Z(n13896) );
  AND U13824 ( .A(n14228), .B(n13745), .Z(n13947) );
  XOR U13825 ( .A(n13967), .B(n13968), .Z(n13893) );
  ANDN U13826 ( .A(n13969), .B(n13970), .Z(n13968) );
  XNOR U13827 ( .A(n13967), .B(n13971), .Z(n13969) );
  XOR U13828 ( .A(n13903), .B(n13972), .Z(n13897) );
  IV U13829 ( .A(n13902), .Z(n13972) );
  XNOR U13830 ( .A(n13899), .B(n13940), .Z(n13902) );
  AND U13831 ( .A(n14441), .B(n13636), .Z(n13940) );
  XOR U13832 ( .A(n13973), .B(n13974), .Z(n13899) );
  ANDN U13833 ( .A(n13975), .B(n13976), .Z(n13974) );
  XNOR U13834 ( .A(n13973), .B(n13977), .Z(n13975) );
  XOR U13835 ( .A(n13909), .B(n13978), .Z(n13903) );
  IV U13836 ( .A(n13908), .Z(n13978) );
  XNOR U13837 ( .A(n13905), .B(n13933), .Z(n13908) );
  AND U13838 ( .A(n14680), .B(n13553), .Z(n13933) );
  XOR U13839 ( .A(n13979), .B(n13980), .Z(n13905) );
  ANDN U13840 ( .A(n13981), .B(n13982), .Z(n13980) );
  XNOR U13841 ( .A(n13979), .B(n13983), .Z(n13981) );
  XOR U13842 ( .A(n13915), .B(n13984), .Z(n13909) );
  IV U13843 ( .A(n13914), .Z(n13984) );
  XNOR U13844 ( .A(n13911), .B(n13926), .Z(n13914) );
  AND U13845 ( .A(n14945), .B(n13496), .Z(n13926) );
  XOR U13846 ( .A(n13985), .B(n13986), .Z(n13911) );
  ANDN U13847 ( .A(n13987), .B(n13988), .Z(n13986) );
  XNOR U13848 ( .A(n13985), .B(n13989), .Z(n13987) );
  XOR U13849 ( .A(n13920), .B(n13990), .Z(n13915) );
  IV U13850 ( .A(n13919), .Z(n13990) );
  XNOR U13851 ( .A(n13916), .B(n13924), .Z(n13919) );
  AND U13852 ( .A(n13470), .B(n15236), .Z(n13924) );
  XOR U13853 ( .A(n13991), .B(n13992), .Z(n13916) );
  ANDN U13854 ( .A(n13993), .B(n13994), .Z(n13992) );
  XNOR U13855 ( .A(n13991), .B(n13995), .Z(n13993) );
  XNOR U13856 ( .A(n13996), .B(n13997), .Z(n13920) );
  ANDN U13857 ( .A(n13998), .B(n13999), .Z(n13997) );
  XNOR U13858 ( .A(n13996), .B(n14000), .Z(n13998) );
  XOR U13859 ( .A(n14001), .B(n14002), .Z(n13921) );
  ANDN U13860 ( .A(n14003), .B(n4652), .Z(n14002) );
  XNOR U13861 ( .A(n14001), .B(n14004), .Z(n4652) );
  XNOR U13862 ( .A(n14001), .B(n4650), .Z(n14003) );
  XOR U13863 ( .A(n13931), .B(n14005), .Z(n4650) );
  IV U13864 ( .A(n13930), .Z(n14005) );
  XNOR U13865 ( .A(n13927), .B(n14006), .Z(n13930) );
  XOR U13866 ( .A(n14007), .B(n14008), .Z(n13927) );
  ANDN U13867 ( .A(n14009), .B(n14010), .Z(n14008) );
  XNOR U13868 ( .A(n14007), .B(n14011), .Z(n14009) );
  XOR U13869 ( .A(n13938), .B(n14012), .Z(n13931) );
  IV U13870 ( .A(n13937), .Z(n14012) );
  XNOR U13871 ( .A(n13934), .B(n14013), .Z(n13937) );
  XOR U13872 ( .A(n14014), .B(n14015), .Z(n13934) );
  ANDN U13873 ( .A(n14016), .B(n14017), .Z(n14015) );
  XNOR U13874 ( .A(n14014), .B(n14018), .Z(n14016) );
  XOR U13875 ( .A(n13945), .B(n14019), .Z(n13938) );
  IV U13876 ( .A(n13944), .Z(n14019) );
  XNOR U13877 ( .A(n13941), .B(n14020), .Z(n13944) );
  XOR U13878 ( .A(n14021), .B(n14022), .Z(n13941) );
  ANDN U13879 ( .A(n14023), .B(n14024), .Z(n14022) );
  XNOR U13880 ( .A(n14021), .B(n14025), .Z(n14023) );
  XOR U13881 ( .A(n13952), .B(n14026), .Z(n13945) );
  IV U13882 ( .A(n13951), .Z(n14026) );
  XNOR U13883 ( .A(n13948), .B(n14027), .Z(n13951) );
  XOR U13884 ( .A(n14028), .B(n14029), .Z(n13948) );
  ANDN U13885 ( .A(n14030), .B(n14031), .Z(n14029) );
  XNOR U13886 ( .A(n14028), .B(n14032), .Z(n14030) );
  XOR U13887 ( .A(n13959), .B(n14033), .Z(n13952) );
  IV U13888 ( .A(n13958), .Z(n14033) );
  XNOR U13889 ( .A(n13955), .B(n14034), .Z(n13958) );
  XOR U13890 ( .A(n14035), .B(n14036), .Z(n13955) );
  ANDN U13891 ( .A(n14037), .B(n14038), .Z(n14036) );
  XNOR U13892 ( .A(n14035), .B(n14039), .Z(n14037) );
  XOR U13893 ( .A(n13965), .B(n14040), .Z(n13959) );
  IV U13894 ( .A(n13964), .Z(n14040) );
  XNOR U13895 ( .A(n13961), .B(n14041), .Z(n13964) );
  XOR U13896 ( .A(n14042), .B(n14043), .Z(n13961) );
  ANDN U13897 ( .A(n14044), .B(n14045), .Z(n14043) );
  XNOR U13898 ( .A(n14042), .B(n14046), .Z(n14044) );
  XOR U13899 ( .A(n13971), .B(n14047), .Z(n13965) );
  IV U13900 ( .A(n13970), .Z(n14047) );
  XNOR U13901 ( .A(n13967), .B(n14034), .Z(n13970) );
  AND U13902 ( .A(n14228), .B(n13880), .Z(n14034) );
  XOR U13903 ( .A(n14048), .B(n14049), .Z(n13967) );
  ANDN U13904 ( .A(n14050), .B(n14051), .Z(n14049) );
  XNOR U13905 ( .A(n14048), .B(n14052), .Z(n14050) );
  XOR U13906 ( .A(n13977), .B(n14053), .Z(n13971) );
  IV U13907 ( .A(n13976), .Z(n14053) );
  XNOR U13908 ( .A(n13973), .B(n14027), .Z(n13976) );
  AND U13909 ( .A(n14441), .B(n13745), .Z(n14027) );
  XOR U13910 ( .A(n14054), .B(n14055), .Z(n13973) );
  ANDN U13911 ( .A(n14056), .B(n14057), .Z(n14055) );
  XNOR U13912 ( .A(n14054), .B(n14058), .Z(n14056) );
  XOR U13913 ( .A(n13983), .B(n14059), .Z(n13977) );
  IV U13914 ( .A(n13982), .Z(n14059) );
  XNOR U13915 ( .A(n13979), .B(n14020), .Z(n13982) );
  AND U13916 ( .A(n14680), .B(n13636), .Z(n14020) );
  XOR U13917 ( .A(n14060), .B(n14061), .Z(n13979) );
  ANDN U13918 ( .A(n14062), .B(n14063), .Z(n14061) );
  XNOR U13919 ( .A(n14060), .B(n14064), .Z(n14062) );
  XOR U13920 ( .A(n13989), .B(n14065), .Z(n13983) );
  IV U13921 ( .A(n13988), .Z(n14065) );
  XNOR U13922 ( .A(n13985), .B(n14013), .Z(n13988) );
  AND U13923 ( .A(n14945), .B(n13553), .Z(n14013) );
  XOR U13924 ( .A(n14066), .B(n14067), .Z(n13985) );
  ANDN U13925 ( .A(n14068), .B(n14069), .Z(n14067) );
  XNOR U13926 ( .A(n14066), .B(n14070), .Z(n14068) );
  XOR U13927 ( .A(n13995), .B(n14071), .Z(n13989) );
  IV U13928 ( .A(n13994), .Z(n14071) );
  XNOR U13929 ( .A(n13991), .B(n14006), .Z(n13994) );
  AND U13930 ( .A(n15236), .B(n13496), .Z(n14006) );
  XOR U13931 ( .A(n14072), .B(n14073), .Z(n13991) );
  ANDN U13932 ( .A(n14074), .B(n14075), .Z(n14073) );
  XNOR U13933 ( .A(n14072), .B(n14076), .Z(n14074) );
  XOR U13934 ( .A(n14000), .B(n14077), .Z(n13995) );
  IV U13935 ( .A(n13999), .Z(n14077) );
  XNOR U13936 ( .A(n13996), .B(n14004), .Z(n13999) );
  AND U13937 ( .A(n13470), .B(n15553), .Z(n14004) );
  XOR U13938 ( .A(n14078), .B(n14079), .Z(n13996) );
  ANDN U13939 ( .A(n14080), .B(n14081), .Z(n14079) );
  XNOR U13940 ( .A(n14078), .B(n14082), .Z(n14080) );
  XNOR U13941 ( .A(n14083), .B(n14084), .Z(n14000) );
  ANDN U13942 ( .A(n14085), .B(n14086), .Z(n14084) );
  XNOR U13943 ( .A(n14083), .B(n14087), .Z(n14085) );
  XOR U13944 ( .A(n14088), .B(n14089), .Z(n14001) );
  ANDN U13945 ( .A(n14090), .B(n4904), .Z(n14089) );
  XNOR U13946 ( .A(n14088), .B(n14091), .Z(n4904) );
  XNOR U13947 ( .A(n14088), .B(n4902), .Z(n14090) );
  XOR U13948 ( .A(n14011), .B(n14092), .Z(n4902) );
  IV U13949 ( .A(n14010), .Z(n14092) );
  XNOR U13950 ( .A(n14007), .B(n14093), .Z(n14010) );
  XOR U13951 ( .A(n14094), .B(n14095), .Z(n14007) );
  ANDN U13952 ( .A(n14096), .B(n14097), .Z(n14095) );
  XNOR U13953 ( .A(n14094), .B(n14098), .Z(n14096) );
  XOR U13954 ( .A(n14018), .B(n14099), .Z(n14011) );
  IV U13955 ( .A(n14017), .Z(n14099) );
  XNOR U13956 ( .A(n14014), .B(n14100), .Z(n14017) );
  XOR U13957 ( .A(n14101), .B(n14102), .Z(n14014) );
  ANDN U13958 ( .A(n14103), .B(n14104), .Z(n14102) );
  XNOR U13959 ( .A(n14101), .B(n14105), .Z(n14103) );
  XOR U13960 ( .A(n14025), .B(n14106), .Z(n14018) );
  IV U13961 ( .A(n14024), .Z(n14106) );
  XNOR U13962 ( .A(n14021), .B(n14107), .Z(n14024) );
  XOR U13963 ( .A(n14108), .B(n14109), .Z(n14021) );
  ANDN U13964 ( .A(n14110), .B(n14111), .Z(n14109) );
  XNOR U13965 ( .A(n14108), .B(n14112), .Z(n14110) );
  XOR U13966 ( .A(n14032), .B(n14113), .Z(n14025) );
  IV U13967 ( .A(n14031), .Z(n14113) );
  XNOR U13968 ( .A(n14028), .B(n14114), .Z(n14031) );
  XOR U13969 ( .A(n14115), .B(n14116), .Z(n14028) );
  ANDN U13970 ( .A(n14117), .B(n14118), .Z(n14116) );
  XNOR U13971 ( .A(n14115), .B(n14119), .Z(n14117) );
  XOR U13972 ( .A(n14039), .B(n14120), .Z(n14032) );
  IV U13973 ( .A(n14038), .Z(n14120) );
  XNOR U13974 ( .A(n14035), .B(n14121), .Z(n14038) );
  XOR U13975 ( .A(n14122), .B(n14123), .Z(n14035) );
  ANDN U13976 ( .A(n14124), .B(n14125), .Z(n14123) );
  XNOR U13977 ( .A(n14122), .B(n14126), .Z(n14124) );
  XOR U13978 ( .A(n14046), .B(n14127), .Z(n14039) );
  IV U13979 ( .A(n14045), .Z(n14127) );
  XNOR U13980 ( .A(n14042), .B(n14128), .Z(n14045) );
  XOR U13981 ( .A(n14129), .B(n14130), .Z(n14042) );
  ANDN U13982 ( .A(n14131), .B(n14132), .Z(n14130) );
  XNOR U13983 ( .A(n14129), .B(n14133), .Z(n14131) );
  XOR U13984 ( .A(n14052), .B(n14134), .Z(n14046) );
  IV U13985 ( .A(n14051), .Z(n14134) );
  XNOR U13986 ( .A(n14048), .B(n14128), .Z(n14051) );
  AND U13987 ( .A(n14228), .B(n14041), .Z(n14128) );
  XOR U13988 ( .A(n14135), .B(n14136), .Z(n14048) );
  ANDN U13989 ( .A(n14137), .B(n14138), .Z(n14136) );
  XNOR U13990 ( .A(n14135), .B(n14139), .Z(n14137) );
  XOR U13991 ( .A(n14058), .B(n14140), .Z(n14052) );
  IV U13992 ( .A(n14057), .Z(n14140) );
  XNOR U13993 ( .A(n14054), .B(n14121), .Z(n14057) );
  AND U13994 ( .A(n14441), .B(n13880), .Z(n14121) );
  XOR U13995 ( .A(n14141), .B(n14142), .Z(n14054) );
  ANDN U13996 ( .A(n14143), .B(n14144), .Z(n14142) );
  XNOR U13997 ( .A(n14141), .B(n14145), .Z(n14143) );
  XOR U13998 ( .A(n14064), .B(n14146), .Z(n14058) );
  IV U13999 ( .A(n14063), .Z(n14146) );
  XNOR U14000 ( .A(n14060), .B(n14114), .Z(n14063) );
  AND U14001 ( .A(n14680), .B(n13745), .Z(n14114) );
  XOR U14002 ( .A(n14147), .B(n14148), .Z(n14060) );
  ANDN U14003 ( .A(n14149), .B(n14150), .Z(n14148) );
  XNOR U14004 ( .A(n14147), .B(n14151), .Z(n14149) );
  XOR U14005 ( .A(n14070), .B(n14152), .Z(n14064) );
  IV U14006 ( .A(n14069), .Z(n14152) );
  XNOR U14007 ( .A(n14066), .B(n14107), .Z(n14069) );
  AND U14008 ( .A(n14945), .B(n13636), .Z(n14107) );
  XOR U14009 ( .A(n14153), .B(n14154), .Z(n14066) );
  ANDN U14010 ( .A(n14155), .B(n14156), .Z(n14154) );
  XNOR U14011 ( .A(n14153), .B(n14157), .Z(n14155) );
  XOR U14012 ( .A(n14076), .B(n14158), .Z(n14070) );
  IV U14013 ( .A(n14075), .Z(n14158) );
  XNOR U14014 ( .A(n14072), .B(n14100), .Z(n14075) );
  AND U14015 ( .A(n15236), .B(n13553), .Z(n14100) );
  XOR U14016 ( .A(n14159), .B(n14160), .Z(n14072) );
  ANDN U14017 ( .A(n14161), .B(n14162), .Z(n14160) );
  XNOR U14018 ( .A(n14159), .B(n14163), .Z(n14161) );
  XOR U14019 ( .A(n14082), .B(n14164), .Z(n14076) );
  IV U14020 ( .A(n14081), .Z(n14164) );
  XNOR U14021 ( .A(n14078), .B(n14093), .Z(n14081) );
  AND U14022 ( .A(n15553), .B(n13496), .Z(n14093) );
  XOR U14023 ( .A(n14165), .B(n14166), .Z(n14078) );
  ANDN U14024 ( .A(n14167), .B(n14168), .Z(n14166) );
  XNOR U14025 ( .A(n14165), .B(n14169), .Z(n14167) );
  XOR U14026 ( .A(n14087), .B(n14170), .Z(n14082) );
  IV U14027 ( .A(n14086), .Z(n14170) );
  XNOR U14028 ( .A(n14083), .B(n14091), .Z(n14086) );
  AND U14029 ( .A(n13470), .B(n15896), .Z(n14091) );
  XOR U14030 ( .A(n14171), .B(n14172), .Z(n14083) );
  ANDN U14031 ( .A(n14173), .B(n14174), .Z(n14172) );
  XNOR U14032 ( .A(n14171), .B(n14175), .Z(n14173) );
  XNOR U14033 ( .A(n14176), .B(n14177), .Z(n14087) );
  ANDN U14034 ( .A(n14178), .B(n14179), .Z(n14177) );
  XNOR U14035 ( .A(n14176), .B(n14180), .Z(n14178) );
  XOR U14036 ( .A(n14181), .B(n14182), .Z(n14088) );
  ANDN U14037 ( .A(n14183), .B(n5163), .Z(n14182) );
  XNOR U14038 ( .A(n14181), .B(n14184), .Z(n5163) );
  XNOR U14039 ( .A(n14181), .B(n5161), .Z(n14183) );
  XOR U14040 ( .A(n14098), .B(n14185), .Z(n5161) );
  IV U14041 ( .A(n14097), .Z(n14185) );
  XNOR U14042 ( .A(n14094), .B(n14186), .Z(n14097) );
  XOR U14043 ( .A(n14187), .B(n14188), .Z(n14094) );
  ANDN U14044 ( .A(n14189), .B(n14190), .Z(n14188) );
  XNOR U14045 ( .A(n14187), .B(n14191), .Z(n14189) );
  XOR U14046 ( .A(n14105), .B(n14192), .Z(n14098) );
  IV U14047 ( .A(n14104), .Z(n14192) );
  XNOR U14048 ( .A(n14101), .B(n14193), .Z(n14104) );
  XOR U14049 ( .A(n14194), .B(n14195), .Z(n14101) );
  ANDN U14050 ( .A(n14196), .B(n14197), .Z(n14195) );
  XNOR U14051 ( .A(n14194), .B(n14198), .Z(n14196) );
  XOR U14052 ( .A(n14112), .B(n14199), .Z(n14105) );
  IV U14053 ( .A(n14111), .Z(n14199) );
  XNOR U14054 ( .A(n14108), .B(n14200), .Z(n14111) );
  XOR U14055 ( .A(n14201), .B(n14202), .Z(n14108) );
  ANDN U14056 ( .A(n14203), .B(n14204), .Z(n14202) );
  XNOR U14057 ( .A(n14201), .B(n14205), .Z(n14203) );
  XOR U14058 ( .A(n14119), .B(n14206), .Z(n14112) );
  IV U14059 ( .A(n14118), .Z(n14206) );
  XNOR U14060 ( .A(n14115), .B(n14207), .Z(n14118) );
  XOR U14061 ( .A(n14208), .B(n14209), .Z(n14115) );
  ANDN U14062 ( .A(n14210), .B(n14211), .Z(n14209) );
  XNOR U14063 ( .A(n14208), .B(n14212), .Z(n14210) );
  XOR U14064 ( .A(n14126), .B(n14213), .Z(n14119) );
  IV U14065 ( .A(n14125), .Z(n14213) );
  XNOR U14066 ( .A(n14122), .B(n14214), .Z(n14125) );
  XOR U14067 ( .A(n14215), .B(n14216), .Z(n14122) );
  ANDN U14068 ( .A(n14217), .B(n14218), .Z(n14216) );
  XNOR U14069 ( .A(n14215), .B(n14219), .Z(n14217) );
  XOR U14070 ( .A(n14133), .B(n14220), .Z(n14126) );
  IV U14071 ( .A(n14132), .Z(n14220) );
  XNOR U14072 ( .A(n14129), .B(n14221), .Z(n14132) );
  XOR U14073 ( .A(n14222), .B(n14223), .Z(n14129) );
  ANDN U14074 ( .A(n14224), .B(n14225), .Z(n14223) );
  XNOR U14075 ( .A(n14222), .B(n14226), .Z(n14224) );
  XOR U14076 ( .A(n14139), .B(n14227), .Z(n14133) );
  IV U14077 ( .A(n14138), .Z(n14227) );
  XNOR U14078 ( .A(n14135), .B(n14228), .Z(n14138) );
  XOR U14079 ( .A(n14229), .B(n14230), .Z(n14135) );
  ANDN U14080 ( .A(n14231), .B(n14232), .Z(n14230) );
  XNOR U14081 ( .A(n14229), .B(n14233), .Z(n14231) );
  XOR U14082 ( .A(n14145), .B(n14234), .Z(n14139) );
  IV U14083 ( .A(n14144), .Z(n14234) );
  XNOR U14084 ( .A(n14141), .B(n14221), .Z(n14144) );
  AND U14085 ( .A(n14441), .B(n14041), .Z(n14221) );
  XOR U14086 ( .A(n14235), .B(n14236), .Z(n14141) );
  ANDN U14087 ( .A(n14237), .B(n14238), .Z(n14236) );
  XNOR U14088 ( .A(n14235), .B(n14239), .Z(n14237) );
  XOR U14089 ( .A(n14151), .B(n14240), .Z(n14145) );
  IV U14090 ( .A(n14150), .Z(n14240) );
  XNOR U14091 ( .A(n14147), .B(n14214), .Z(n14150) );
  AND U14092 ( .A(n14680), .B(n13880), .Z(n14214) );
  XOR U14093 ( .A(n14241), .B(n14242), .Z(n14147) );
  ANDN U14094 ( .A(n14243), .B(n14244), .Z(n14242) );
  XNOR U14095 ( .A(n14241), .B(n14245), .Z(n14243) );
  XOR U14096 ( .A(n14157), .B(n14246), .Z(n14151) );
  IV U14097 ( .A(n14156), .Z(n14246) );
  XNOR U14098 ( .A(n14153), .B(n14207), .Z(n14156) );
  AND U14099 ( .A(n14945), .B(n13745), .Z(n14207) );
  XOR U14100 ( .A(n14247), .B(n14248), .Z(n14153) );
  ANDN U14101 ( .A(n14249), .B(n14250), .Z(n14248) );
  XNOR U14102 ( .A(n14247), .B(n14251), .Z(n14249) );
  XOR U14103 ( .A(n14163), .B(n14252), .Z(n14157) );
  IV U14104 ( .A(n14162), .Z(n14252) );
  XNOR U14105 ( .A(n14159), .B(n14200), .Z(n14162) );
  AND U14106 ( .A(n15236), .B(n13636), .Z(n14200) );
  XOR U14107 ( .A(n14253), .B(n14254), .Z(n14159) );
  ANDN U14108 ( .A(n14255), .B(n14256), .Z(n14254) );
  XNOR U14109 ( .A(n14253), .B(n14257), .Z(n14255) );
  XOR U14110 ( .A(n14169), .B(n14258), .Z(n14163) );
  IV U14111 ( .A(n14168), .Z(n14258) );
  XNOR U14112 ( .A(n14165), .B(n14193), .Z(n14168) );
  AND U14113 ( .A(n15553), .B(n13553), .Z(n14193) );
  XOR U14114 ( .A(n14259), .B(n14260), .Z(n14165) );
  ANDN U14115 ( .A(n14261), .B(n14262), .Z(n14260) );
  XNOR U14116 ( .A(n14259), .B(n14263), .Z(n14261) );
  XOR U14117 ( .A(n14175), .B(n14264), .Z(n14169) );
  IV U14118 ( .A(n14174), .Z(n14264) );
  XNOR U14119 ( .A(n14171), .B(n14186), .Z(n14174) );
  AND U14120 ( .A(n15896), .B(n13496), .Z(n14186) );
  XOR U14121 ( .A(n14265), .B(n14266), .Z(n14171) );
  ANDN U14122 ( .A(n14267), .B(n14268), .Z(n14266) );
  XNOR U14123 ( .A(n14265), .B(n14269), .Z(n14267) );
  XOR U14124 ( .A(n14180), .B(n14270), .Z(n14175) );
  IV U14125 ( .A(n14179), .Z(n14270) );
  XNOR U14126 ( .A(n14176), .B(n14184), .Z(n14179) );
  AND U14127 ( .A(n13470), .B(n16265), .Z(n14184) );
  XOR U14128 ( .A(n14271), .B(n14272), .Z(n14176) );
  ANDN U14129 ( .A(n14273), .B(n14274), .Z(n14272) );
  XNOR U14130 ( .A(n14271), .B(n14275), .Z(n14273) );
  XNOR U14131 ( .A(n14276), .B(n14277), .Z(n14180) );
  ANDN U14132 ( .A(n14278), .B(n14279), .Z(n14277) );
  XNOR U14133 ( .A(n14276), .B(n14280), .Z(n14278) );
  XOR U14134 ( .A(n14281), .B(n14282), .Z(n14181) );
  ANDN U14135 ( .A(n14283), .B(n5428), .Z(n14282) );
  XNOR U14136 ( .A(n14281), .B(n14284), .Z(n5428) );
  XNOR U14137 ( .A(n14281), .B(n5426), .Z(n14283) );
  XOR U14138 ( .A(n14191), .B(n14285), .Z(n5426) );
  IV U14139 ( .A(n14190), .Z(n14285) );
  XNOR U14140 ( .A(n14187), .B(n14286), .Z(n14190) );
  XOR U14141 ( .A(n14287), .B(n14288), .Z(n14187) );
  ANDN U14142 ( .A(n14289), .B(n14290), .Z(n14288) );
  XNOR U14143 ( .A(n14287), .B(n14291), .Z(n14289) );
  XOR U14144 ( .A(n14198), .B(n14292), .Z(n14191) );
  IV U14145 ( .A(n14197), .Z(n14292) );
  XNOR U14146 ( .A(n14194), .B(n14293), .Z(n14197) );
  XOR U14147 ( .A(n14294), .B(n14295), .Z(n14194) );
  ANDN U14148 ( .A(n14296), .B(n14297), .Z(n14295) );
  XNOR U14149 ( .A(n14294), .B(n14298), .Z(n14296) );
  XOR U14150 ( .A(n14205), .B(n14299), .Z(n14198) );
  IV U14151 ( .A(n14204), .Z(n14299) );
  XNOR U14152 ( .A(n14201), .B(n14300), .Z(n14204) );
  XOR U14153 ( .A(n14301), .B(n14302), .Z(n14201) );
  ANDN U14154 ( .A(n14303), .B(n14304), .Z(n14302) );
  XNOR U14155 ( .A(n14301), .B(n14305), .Z(n14303) );
  XOR U14156 ( .A(n14212), .B(n14306), .Z(n14205) );
  IV U14157 ( .A(n14211), .Z(n14306) );
  XNOR U14158 ( .A(n14208), .B(n14307), .Z(n14211) );
  XOR U14159 ( .A(n14308), .B(n14309), .Z(n14208) );
  ANDN U14160 ( .A(n14310), .B(n14311), .Z(n14309) );
  XNOR U14161 ( .A(n14308), .B(n14312), .Z(n14310) );
  XOR U14162 ( .A(n14219), .B(n14313), .Z(n14212) );
  IV U14163 ( .A(n14218), .Z(n14313) );
  XNOR U14164 ( .A(n14215), .B(n14314), .Z(n14218) );
  XOR U14165 ( .A(n14315), .B(n14316), .Z(n14215) );
  ANDN U14166 ( .A(n14317), .B(n14318), .Z(n14316) );
  XNOR U14167 ( .A(n14315), .B(n14319), .Z(n14317) );
  XOR U14168 ( .A(n14226), .B(n14320), .Z(n14219) );
  IV U14169 ( .A(n14225), .Z(n14320) );
  XNOR U14170 ( .A(n14222), .B(n14321), .Z(n14225) );
  XOR U14171 ( .A(n14322), .B(n14323), .Z(n14222) );
  ANDN U14172 ( .A(n14324), .B(n14325), .Z(n14323) );
  XNOR U14173 ( .A(n14322), .B(n14326), .Z(n14324) );
  XOR U14174 ( .A(n14233), .B(n14327), .Z(n14226) );
  IV U14175 ( .A(n14232), .Z(n14327) );
  XNOR U14176 ( .A(n14229), .B(n14328), .Z(n14232) );
  XOR U14177 ( .A(n14329), .B(n14330), .Z(n14229) );
  ANDN U14178 ( .A(n14331), .B(n14332), .Z(n14330) );
  XNOR U14179 ( .A(n14329), .B(n14333), .Z(n14331) );
  XOR U14180 ( .A(n14239), .B(n14334), .Z(n14233) );
  IV U14181 ( .A(n14238), .Z(n14334) );
  XNOR U14182 ( .A(n14235), .B(n14328), .Z(n14238) );
  AND U14183 ( .A(n14441), .B(n14228), .Z(n14328) );
  XOR U14184 ( .A(n14335), .B(n14336), .Z(n14235) );
  ANDN U14185 ( .A(n14337), .B(n14338), .Z(n14336) );
  XNOR U14186 ( .A(n14335), .B(n14339), .Z(n14337) );
  XOR U14187 ( .A(n14245), .B(n14340), .Z(n14239) );
  IV U14188 ( .A(n14244), .Z(n14340) );
  XNOR U14189 ( .A(n14241), .B(n14321), .Z(n14244) );
  AND U14190 ( .A(n14680), .B(n14041), .Z(n14321) );
  XOR U14191 ( .A(n14341), .B(n14342), .Z(n14241) );
  ANDN U14192 ( .A(n14343), .B(n14344), .Z(n14342) );
  XNOR U14193 ( .A(n14341), .B(n14345), .Z(n14343) );
  XOR U14194 ( .A(n14251), .B(n14346), .Z(n14245) );
  IV U14195 ( .A(n14250), .Z(n14346) );
  XNOR U14196 ( .A(n14247), .B(n14314), .Z(n14250) );
  AND U14197 ( .A(n14945), .B(n13880), .Z(n14314) );
  XOR U14198 ( .A(n14347), .B(n14348), .Z(n14247) );
  ANDN U14199 ( .A(n14349), .B(n14350), .Z(n14348) );
  XNOR U14200 ( .A(n14347), .B(n14351), .Z(n14349) );
  XOR U14201 ( .A(n14257), .B(n14352), .Z(n14251) );
  IV U14202 ( .A(n14256), .Z(n14352) );
  XNOR U14203 ( .A(n14253), .B(n14307), .Z(n14256) );
  AND U14204 ( .A(n15236), .B(n13745), .Z(n14307) );
  XOR U14205 ( .A(n14353), .B(n14354), .Z(n14253) );
  ANDN U14206 ( .A(n14355), .B(n14356), .Z(n14354) );
  XNOR U14207 ( .A(n14353), .B(n14357), .Z(n14355) );
  XOR U14208 ( .A(n14263), .B(n14358), .Z(n14257) );
  IV U14209 ( .A(n14262), .Z(n14358) );
  XNOR U14210 ( .A(n14259), .B(n14300), .Z(n14262) );
  AND U14211 ( .A(n15553), .B(n13636), .Z(n14300) );
  XOR U14212 ( .A(n14359), .B(n14360), .Z(n14259) );
  ANDN U14213 ( .A(n14361), .B(n14362), .Z(n14360) );
  XNOR U14214 ( .A(n14359), .B(n14363), .Z(n14361) );
  XOR U14215 ( .A(n14269), .B(n14364), .Z(n14263) );
  IV U14216 ( .A(n14268), .Z(n14364) );
  XNOR U14217 ( .A(n14265), .B(n14293), .Z(n14268) );
  AND U14218 ( .A(n15896), .B(n13553), .Z(n14293) );
  XOR U14219 ( .A(n14365), .B(n14366), .Z(n14265) );
  ANDN U14220 ( .A(n14367), .B(n14368), .Z(n14366) );
  XNOR U14221 ( .A(n14365), .B(n14369), .Z(n14367) );
  XOR U14222 ( .A(n14275), .B(n14370), .Z(n14269) );
  IV U14223 ( .A(n14274), .Z(n14370) );
  XNOR U14224 ( .A(n14271), .B(n14286), .Z(n14274) );
  AND U14225 ( .A(n16265), .B(n13496), .Z(n14286) );
  XOR U14226 ( .A(n14371), .B(n14372), .Z(n14271) );
  ANDN U14227 ( .A(n14373), .B(n14374), .Z(n14372) );
  XNOR U14228 ( .A(n14371), .B(n14375), .Z(n14373) );
  XOR U14229 ( .A(n14280), .B(n14376), .Z(n14275) );
  IV U14230 ( .A(n14279), .Z(n14376) );
  XNOR U14231 ( .A(n14276), .B(n14284), .Z(n14279) );
  AND U14232 ( .A(n13470), .B(n16657), .Z(n14284) );
  XOR U14233 ( .A(n14377), .B(n14378), .Z(n14276) );
  ANDN U14234 ( .A(n14379), .B(n14380), .Z(n14378) );
  XNOR U14235 ( .A(n14377), .B(n14381), .Z(n14379) );
  XNOR U14236 ( .A(n14382), .B(n14383), .Z(n14280) );
  ANDN U14237 ( .A(n14384), .B(n14385), .Z(n14383) );
  XNOR U14238 ( .A(n14382), .B(n14386), .Z(n14384) );
  XOR U14239 ( .A(n14387), .B(n14388), .Z(n14281) );
  ANDN U14240 ( .A(n14389), .B(n5700), .Z(n14388) );
  XNOR U14241 ( .A(n14387), .B(n14390), .Z(n5700) );
  XNOR U14242 ( .A(n14387), .B(n5698), .Z(n14389) );
  XOR U14243 ( .A(n14291), .B(n14391), .Z(n5698) );
  IV U14244 ( .A(n14290), .Z(n14391) );
  XNOR U14245 ( .A(n14287), .B(n14392), .Z(n14290) );
  XOR U14246 ( .A(n14393), .B(n14394), .Z(n14287) );
  ANDN U14247 ( .A(n14395), .B(n14396), .Z(n14394) );
  XNOR U14248 ( .A(n14393), .B(n14397), .Z(n14395) );
  XOR U14249 ( .A(n14298), .B(n14398), .Z(n14291) );
  IV U14250 ( .A(n14297), .Z(n14398) );
  XNOR U14251 ( .A(n14294), .B(n14399), .Z(n14297) );
  XOR U14252 ( .A(n14400), .B(n14401), .Z(n14294) );
  ANDN U14253 ( .A(n14402), .B(n14403), .Z(n14401) );
  XNOR U14254 ( .A(n14400), .B(n14404), .Z(n14402) );
  XOR U14255 ( .A(n14305), .B(n14405), .Z(n14298) );
  IV U14256 ( .A(n14304), .Z(n14405) );
  XNOR U14257 ( .A(n14301), .B(n14406), .Z(n14304) );
  XOR U14258 ( .A(n14407), .B(n14408), .Z(n14301) );
  ANDN U14259 ( .A(n14409), .B(n14410), .Z(n14408) );
  XNOR U14260 ( .A(n14407), .B(n14411), .Z(n14409) );
  XOR U14261 ( .A(n14312), .B(n14412), .Z(n14305) );
  IV U14262 ( .A(n14311), .Z(n14412) );
  XNOR U14263 ( .A(n14308), .B(n14413), .Z(n14311) );
  XOR U14264 ( .A(n14414), .B(n14415), .Z(n14308) );
  ANDN U14265 ( .A(n14416), .B(n14417), .Z(n14415) );
  XNOR U14266 ( .A(n14414), .B(n14418), .Z(n14416) );
  XOR U14267 ( .A(n14319), .B(n14419), .Z(n14312) );
  IV U14268 ( .A(n14318), .Z(n14419) );
  XNOR U14269 ( .A(n14315), .B(n14420), .Z(n14318) );
  XOR U14270 ( .A(n14421), .B(n14422), .Z(n14315) );
  ANDN U14271 ( .A(n14423), .B(n14424), .Z(n14422) );
  XNOR U14272 ( .A(n14421), .B(n14425), .Z(n14423) );
  XOR U14273 ( .A(n14326), .B(n14426), .Z(n14319) );
  IV U14274 ( .A(n14325), .Z(n14426) );
  XNOR U14275 ( .A(n14322), .B(n14427), .Z(n14325) );
  XOR U14276 ( .A(n14428), .B(n14429), .Z(n14322) );
  ANDN U14277 ( .A(n14430), .B(n14431), .Z(n14429) );
  XNOR U14278 ( .A(n14428), .B(n14432), .Z(n14430) );
  XOR U14279 ( .A(n14333), .B(n14433), .Z(n14326) );
  IV U14280 ( .A(n14332), .Z(n14433) );
  XNOR U14281 ( .A(n14329), .B(n14434), .Z(n14332) );
  XOR U14282 ( .A(n14435), .B(n14436), .Z(n14329) );
  ANDN U14283 ( .A(n14437), .B(n14438), .Z(n14436) );
  XNOR U14284 ( .A(n14435), .B(n14439), .Z(n14437) );
  XOR U14285 ( .A(n14339), .B(n14440), .Z(n14333) );
  IV U14286 ( .A(n14338), .Z(n14440) );
  XNOR U14287 ( .A(n14335), .B(n14441), .Z(n14338) );
  XOR U14288 ( .A(n14442), .B(n14443), .Z(n14335) );
  ANDN U14289 ( .A(n14444), .B(n14445), .Z(n14443) );
  XNOR U14290 ( .A(n14442), .B(n14446), .Z(n14444) );
  XOR U14291 ( .A(n14345), .B(n14447), .Z(n14339) );
  IV U14292 ( .A(n14344), .Z(n14447) );
  XNOR U14293 ( .A(n14341), .B(n14434), .Z(n14344) );
  AND U14294 ( .A(n14680), .B(n14228), .Z(n14434) );
  XOR U14295 ( .A(n14448), .B(n14449), .Z(n14341) );
  ANDN U14296 ( .A(n14450), .B(n14451), .Z(n14449) );
  XNOR U14297 ( .A(n14448), .B(n14452), .Z(n14450) );
  XOR U14298 ( .A(n14351), .B(n14453), .Z(n14345) );
  IV U14299 ( .A(n14350), .Z(n14453) );
  XNOR U14300 ( .A(n14347), .B(n14427), .Z(n14350) );
  AND U14301 ( .A(n14945), .B(n14041), .Z(n14427) );
  XOR U14302 ( .A(n14454), .B(n14455), .Z(n14347) );
  ANDN U14303 ( .A(n14456), .B(n14457), .Z(n14455) );
  XNOR U14304 ( .A(n14454), .B(n14458), .Z(n14456) );
  XOR U14305 ( .A(n14357), .B(n14459), .Z(n14351) );
  IV U14306 ( .A(n14356), .Z(n14459) );
  XNOR U14307 ( .A(n14353), .B(n14420), .Z(n14356) );
  AND U14308 ( .A(n15236), .B(n13880), .Z(n14420) );
  XOR U14309 ( .A(n14460), .B(n14461), .Z(n14353) );
  ANDN U14310 ( .A(n14462), .B(n14463), .Z(n14461) );
  XNOR U14311 ( .A(n14460), .B(n14464), .Z(n14462) );
  XOR U14312 ( .A(n14363), .B(n14465), .Z(n14357) );
  IV U14313 ( .A(n14362), .Z(n14465) );
  XNOR U14314 ( .A(n14359), .B(n14413), .Z(n14362) );
  AND U14315 ( .A(n15553), .B(n13745), .Z(n14413) );
  XOR U14316 ( .A(n14466), .B(n14467), .Z(n14359) );
  ANDN U14317 ( .A(n14468), .B(n14469), .Z(n14467) );
  XNOR U14318 ( .A(n14466), .B(n14470), .Z(n14468) );
  XOR U14319 ( .A(n14369), .B(n14471), .Z(n14363) );
  IV U14320 ( .A(n14368), .Z(n14471) );
  XNOR U14321 ( .A(n14365), .B(n14406), .Z(n14368) );
  AND U14322 ( .A(n15896), .B(n13636), .Z(n14406) );
  XOR U14323 ( .A(n14472), .B(n14473), .Z(n14365) );
  ANDN U14324 ( .A(n14474), .B(n14475), .Z(n14473) );
  XNOR U14325 ( .A(n14472), .B(n14476), .Z(n14474) );
  XOR U14326 ( .A(n14375), .B(n14477), .Z(n14369) );
  IV U14327 ( .A(n14374), .Z(n14477) );
  XNOR U14328 ( .A(n14371), .B(n14399), .Z(n14374) );
  AND U14329 ( .A(n16265), .B(n13553), .Z(n14399) );
  XOR U14330 ( .A(n14478), .B(n14479), .Z(n14371) );
  ANDN U14331 ( .A(n14480), .B(n14481), .Z(n14479) );
  XNOR U14332 ( .A(n14478), .B(n14482), .Z(n14480) );
  XOR U14333 ( .A(n14381), .B(n14483), .Z(n14375) );
  IV U14334 ( .A(n14380), .Z(n14483) );
  XNOR U14335 ( .A(n14377), .B(n14392), .Z(n14380) );
  AND U14336 ( .A(n16657), .B(n13496), .Z(n14392) );
  XOR U14337 ( .A(n14484), .B(n14485), .Z(n14377) );
  ANDN U14338 ( .A(n14486), .B(n14487), .Z(n14485) );
  XNOR U14339 ( .A(n14484), .B(n14488), .Z(n14486) );
  XOR U14340 ( .A(n14386), .B(n14489), .Z(n14381) );
  IV U14341 ( .A(n14385), .Z(n14489) );
  XNOR U14342 ( .A(n14382), .B(n14390), .Z(n14385) );
  AND U14343 ( .A(n13470), .B(n17567), .Z(n14390) );
  XOR U14344 ( .A(n14490), .B(n14491), .Z(n14382) );
  ANDN U14345 ( .A(n14492), .B(n14493), .Z(n14491) );
  XNOR U14346 ( .A(n14490), .B(n14494), .Z(n14492) );
  XNOR U14347 ( .A(n14495), .B(n14496), .Z(n14386) );
  ANDN U14348 ( .A(n14497), .B(n14498), .Z(n14496) );
  XNOR U14349 ( .A(n14495), .B(n14499), .Z(n14497) );
  XOR U14350 ( .A(n14500), .B(n14501), .Z(n14387) );
  ANDN U14351 ( .A(n14502), .B(n5978), .Z(n14501) );
  XNOR U14352 ( .A(n14500), .B(n14503), .Z(n5978) );
  XNOR U14353 ( .A(n14500), .B(n5976), .Z(n14502) );
  XOR U14354 ( .A(n14397), .B(n14504), .Z(n5976) );
  IV U14355 ( .A(n14396), .Z(n14504) );
  XNOR U14356 ( .A(n14393), .B(n14505), .Z(n14396) );
  XOR U14357 ( .A(n14506), .B(n14507), .Z(n14393) );
  ANDN U14358 ( .A(n14508), .B(n14509), .Z(n14507) );
  XNOR U14359 ( .A(n14506), .B(n14510), .Z(n14508) );
  XOR U14360 ( .A(n14404), .B(n14511), .Z(n14397) );
  IV U14361 ( .A(n14403), .Z(n14511) );
  XNOR U14362 ( .A(n14400), .B(n14512), .Z(n14403) );
  XOR U14363 ( .A(n14513), .B(n14514), .Z(n14400) );
  ANDN U14364 ( .A(n14515), .B(n14516), .Z(n14514) );
  XNOR U14365 ( .A(n14513), .B(n14517), .Z(n14515) );
  XOR U14366 ( .A(n14411), .B(n14518), .Z(n14404) );
  IV U14367 ( .A(n14410), .Z(n14518) );
  XNOR U14368 ( .A(n14407), .B(n14519), .Z(n14410) );
  XOR U14369 ( .A(n14520), .B(n14521), .Z(n14407) );
  ANDN U14370 ( .A(n14522), .B(n14523), .Z(n14521) );
  XNOR U14371 ( .A(n14520), .B(n14524), .Z(n14522) );
  XOR U14372 ( .A(n14418), .B(n14525), .Z(n14411) );
  IV U14373 ( .A(n14417), .Z(n14525) );
  XNOR U14374 ( .A(n14414), .B(n14526), .Z(n14417) );
  XOR U14375 ( .A(n14527), .B(n14528), .Z(n14414) );
  ANDN U14376 ( .A(n14529), .B(n14530), .Z(n14528) );
  XNOR U14377 ( .A(n14527), .B(n14531), .Z(n14529) );
  XOR U14378 ( .A(n14425), .B(n14532), .Z(n14418) );
  IV U14379 ( .A(n14424), .Z(n14532) );
  XNOR U14380 ( .A(n14421), .B(n14533), .Z(n14424) );
  XOR U14381 ( .A(n14534), .B(n14535), .Z(n14421) );
  ANDN U14382 ( .A(n14536), .B(n14537), .Z(n14535) );
  XNOR U14383 ( .A(n14534), .B(n14538), .Z(n14536) );
  XOR U14384 ( .A(n14432), .B(n14539), .Z(n14425) );
  IV U14385 ( .A(n14431), .Z(n14539) );
  XNOR U14386 ( .A(n14428), .B(n14540), .Z(n14431) );
  XOR U14387 ( .A(n14541), .B(n14542), .Z(n14428) );
  ANDN U14388 ( .A(n14543), .B(n14544), .Z(n14542) );
  XNOR U14389 ( .A(n14541), .B(n14545), .Z(n14543) );
  XOR U14390 ( .A(n14439), .B(n14546), .Z(n14432) );
  IV U14391 ( .A(n14438), .Z(n14546) );
  XNOR U14392 ( .A(n14435), .B(n14547), .Z(n14438) );
  XOR U14393 ( .A(n14548), .B(n14549), .Z(n14435) );
  ANDN U14394 ( .A(n14550), .B(n14551), .Z(n14549) );
  XNOR U14395 ( .A(n14548), .B(n14552), .Z(n14550) );
  XOR U14396 ( .A(n14446), .B(n14553), .Z(n14439) );
  IV U14397 ( .A(n14445), .Z(n14553) );
  XNOR U14398 ( .A(n14442), .B(n14554), .Z(n14445) );
  XOR U14399 ( .A(n14555), .B(n14556), .Z(n14442) );
  ANDN U14400 ( .A(n14557), .B(n14558), .Z(n14556) );
  XNOR U14401 ( .A(n14555), .B(n14559), .Z(n14557) );
  XOR U14402 ( .A(n14452), .B(n14560), .Z(n14446) );
  IV U14403 ( .A(n14451), .Z(n14560) );
  XNOR U14404 ( .A(n14448), .B(n14554), .Z(n14451) );
  AND U14405 ( .A(n14680), .B(n14441), .Z(n14554) );
  XOR U14406 ( .A(n14561), .B(n14562), .Z(n14448) );
  ANDN U14407 ( .A(n14563), .B(n14564), .Z(n14562) );
  XNOR U14408 ( .A(n14561), .B(n14565), .Z(n14563) );
  XOR U14409 ( .A(n14458), .B(n14566), .Z(n14452) );
  IV U14410 ( .A(n14457), .Z(n14566) );
  XNOR U14411 ( .A(n14454), .B(n14547), .Z(n14457) );
  AND U14412 ( .A(n14945), .B(n14228), .Z(n14547) );
  XOR U14413 ( .A(n14567), .B(n14568), .Z(n14454) );
  ANDN U14414 ( .A(n14569), .B(n14570), .Z(n14568) );
  XNOR U14415 ( .A(n14567), .B(n14571), .Z(n14569) );
  XOR U14416 ( .A(n14464), .B(n14572), .Z(n14458) );
  IV U14417 ( .A(n14463), .Z(n14572) );
  XNOR U14418 ( .A(n14460), .B(n14540), .Z(n14463) );
  AND U14419 ( .A(n15236), .B(n14041), .Z(n14540) );
  XOR U14420 ( .A(n14573), .B(n14574), .Z(n14460) );
  ANDN U14421 ( .A(n14575), .B(n14576), .Z(n14574) );
  XNOR U14422 ( .A(n14573), .B(n14577), .Z(n14575) );
  XOR U14423 ( .A(n14470), .B(n14578), .Z(n14464) );
  IV U14424 ( .A(n14469), .Z(n14578) );
  XNOR U14425 ( .A(n14466), .B(n14533), .Z(n14469) );
  AND U14426 ( .A(n15553), .B(n13880), .Z(n14533) );
  XOR U14427 ( .A(n14579), .B(n14580), .Z(n14466) );
  ANDN U14428 ( .A(n14581), .B(n14582), .Z(n14580) );
  XNOR U14429 ( .A(n14579), .B(n14583), .Z(n14581) );
  XOR U14430 ( .A(n14476), .B(n14584), .Z(n14470) );
  IV U14431 ( .A(n14475), .Z(n14584) );
  XNOR U14432 ( .A(n14472), .B(n14526), .Z(n14475) );
  AND U14433 ( .A(n15896), .B(n13745), .Z(n14526) );
  XOR U14434 ( .A(n14585), .B(n14586), .Z(n14472) );
  ANDN U14435 ( .A(n14587), .B(n14588), .Z(n14586) );
  XNOR U14436 ( .A(n14585), .B(n14589), .Z(n14587) );
  XOR U14437 ( .A(n14482), .B(n14590), .Z(n14476) );
  IV U14438 ( .A(n14481), .Z(n14590) );
  XNOR U14439 ( .A(n14478), .B(n14519), .Z(n14481) );
  AND U14440 ( .A(n16265), .B(n13636), .Z(n14519) );
  XOR U14441 ( .A(n14591), .B(n14592), .Z(n14478) );
  ANDN U14442 ( .A(n14593), .B(n14594), .Z(n14592) );
  XNOR U14443 ( .A(n14591), .B(n14595), .Z(n14593) );
  XOR U14444 ( .A(n14488), .B(n14596), .Z(n14482) );
  IV U14445 ( .A(n14487), .Z(n14596) );
  XNOR U14446 ( .A(n14484), .B(n14512), .Z(n14487) );
  AND U14447 ( .A(n16657), .B(n13553), .Z(n14512) );
  XOR U14448 ( .A(n14597), .B(n14598), .Z(n14484) );
  ANDN U14449 ( .A(n14599), .B(n14600), .Z(n14598) );
  XNOR U14450 ( .A(n14597), .B(n14601), .Z(n14599) );
  XOR U14451 ( .A(n14494), .B(n14602), .Z(n14488) );
  IV U14452 ( .A(n14493), .Z(n14602) );
  XNOR U14453 ( .A(n14490), .B(n14505), .Z(n14493) );
  AND U14454 ( .A(n17567), .B(n13496), .Z(n14505) );
  XOR U14455 ( .A(n14603), .B(n14604), .Z(n14490) );
  ANDN U14456 ( .A(n14605), .B(n14606), .Z(n14604) );
  XNOR U14457 ( .A(n14603), .B(n14607), .Z(n14605) );
  XOR U14458 ( .A(n14499), .B(n14608), .Z(n14494) );
  IV U14459 ( .A(n14498), .Z(n14608) );
  XNOR U14460 ( .A(n14495), .B(n14503), .Z(n14498) );
  AND U14461 ( .A(n13470), .B(n17688), .Z(n14503) );
  XOR U14462 ( .A(n14609), .B(n14610), .Z(n14495) );
  ANDN U14463 ( .A(n14611), .B(n14612), .Z(n14610) );
  XNOR U14464 ( .A(n14609), .B(n14613), .Z(n14611) );
  XNOR U14465 ( .A(n14614), .B(n14615), .Z(n14499) );
  ANDN U14466 ( .A(n14616), .B(n14617), .Z(n14615) );
  XNOR U14467 ( .A(n14614), .B(n14618), .Z(n14616) );
  XOR U14468 ( .A(n14619), .B(n14620), .Z(n14500) );
  ANDN U14469 ( .A(n14621), .B(n6261), .Z(n14620) );
  XNOR U14470 ( .A(n14619), .B(n14622), .Z(n6261) );
  XNOR U14471 ( .A(n14619), .B(n6259), .Z(n14621) );
  XOR U14472 ( .A(n14510), .B(n14623), .Z(n6259) );
  IV U14473 ( .A(n14509), .Z(n14623) );
  XNOR U14474 ( .A(n14506), .B(n14624), .Z(n14509) );
  XOR U14475 ( .A(n14625), .B(n14626), .Z(n14506) );
  ANDN U14476 ( .A(n14627), .B(n14628), .Z(n14626) );
  XNOR U14477 ( .A(n14625), .B(n14629), .Z(n14627) );
  XOR U14478 ( .A(n14517), .B(n14630), .Z(n14510) );
  IV U14479 ( .A(n14516), .Z(n14630) );
  XNOR U14480 ( .A(n14513), .B(n14631), .Z(n14516) );
  XOR U14481 ( .A(n14632), .B(n14633), .Z(n14513) );
  ANDN U14482 ( .A(n14634), .B(n14635), .Z(n14633) );
  XNOR U14483 ( .A(n14632), .B(n14636), .Z(n14634) );
  XOR U14484 ( .A(n14524), .B(n14637), .Z(n14517) );
  IV U14485 ( .A(n14523), .Z(n14637) );
  XNOR U14486 ( .A(n14520), .B(n14638), .Z(n14523) );
  XOR U14487 ( .A(n14639), .B(n14640), .Z(n14520) );
  ANDN U14488 ( .A(n14641), .B(n14642), .Z(n14640) );
  XNOR U14489 ( .A(n14639), .B(n14643), .Z(n14641) );
  XOR U14490 ( .A(n14531), .B(n14644), .Z(n14524) );
  IV U14491 ( .A(n14530), .Z(n14644) );
  XNOR U14492 ( .A(n14527), .B(n14645), .Z(n14530) );
  XOR U14493 ( .A(n14646), .B(n14647), .Z(n14527) );
  ANDN U14494 ( .A(n14648), .B(n14649), .Z(n14647) );
  XNOR U14495 ( .A(n14646), .B(n14650), .Z(n14648) );
  XOR U14496 ( .A(n14538), .B(n14651), .Z(n14531) );
  IV U14497 ( .A(n14537), .Z(n14651) );
  XNOR U14498 ( .A(n14534), .B(n14652), .Z(n14537) );
  XOR U14499 ( .A(n14653), .B(n14654), .Z(n14534) );
  ANDN U14500 ( .A(n14655), .B(n14656), .Z(n14654) );
  XNOR U14501 ( .A(n14653), .B(n14657), .Z(n14655) );
  XOR U14502 ( .A(n14545), .B(n14658), .Z(n14538) );
  IV U14503 ( .A(n14544), .Z(n14658) );
  XNOR U14504 ( .A(n14541), .B(n14659), .Z(n14544) );
  XOR U14505 ( .A(n14660), .B(n14661), .Z(n14541) );
  ANDN U14506 ( .A(n14662), .B(n14663), .Z(n14661) );
  XNOR U14507 ( .A(n14660), .B(n14664), .Z(n14662) );
  XOR U14508 ( .A(n14552), .B(n14665), .Z(n14545) );
  IV U14509 ( .A(n14551), .Z(n14665) );
  XNOR U14510 ( .A(n14548), .B(n14666), .Z(n14551) );
  XOR U14511 ( .A(n14667), .B(n14668), .Z(n14548) );
  ANDN U14512 ( .A(n14669), .B(n14670), .Z(n14668) );
  XNOR U14513 ( .A(n14667), .B(n14671), .Z(n14669) );
  XOR U14514 ( .A(n14559), .B(n14672), .Z(n14552) );
  IV U14515 ( .A(n14558), .Z(n14672) );
  XNOR U14516 ( .A(n14555), .B(n14673), .Z(n14558) );
  XOR U14517 ( .A(n14674), .B(n14675), .Z(n14555) );
  ANDN U14518 ( .A(n14676), .B(n14677), .Z(n14675) );
  XNOR U14519 ( .A(n14674), .B(n14678), .Z(n14676) );
  XOR U14520 ( .A(n14565), .B(n14679), .Z(n14559) );
  IV U14521 ( .A(n14564), .Z(n14679) );
  XNOR U14522 ( .A(n14561), .B(n14680), .Z(n14564) );
  XOR U14523 ( .A(n14681), .B(n14682), .Z(n14561) );
  ANDN U14524 ( .A(n14683), .B(n14684), .Z(n14682) );
  XNOR U14525 ( .A(n14681), .B(n14685), .Z(n14683) );
  XOR U14526 ( .A(n14571), .B(n14686), .Z(n14565) );
  IV U14527 ( .A(n14570), .Z(n14686) );
  XNOR U14528 ( .A(n14567), .B(n14673), .Z(n14570) );
  AND U14529 ( .A(n14945), .B(n14441), .Z(n14673) );
  XOR U14530 ( .A(n14687), .B(n14688), .Z(n14567) );
  ANDN U14531 ( .A(n14689), .B(n14690), .Z(n14688) );
  XNOR U14532 ( .A(n14687), .B(n14691), .Z(n14689) );
  XOR U14533 ( .A(n14577), .B(n14692), .Z(n14571) );
  IV U14534 ( .A(n14576), .Z(n14692) );
  XNOR U14535 ( .A(n14573), .B(n14666), .Z(n14576) );
  AND U14536 ( .A(n15236), .B(n14228), .Z(n14666) );
  XOR U14537 ( .A(n14693), .B(n14694), .Z(n14573) );
  ANDN U14538 ( .A(n14695), .B(n14696), .Z(n14694) );
  XNOR U14539 ( .A(n14693), .B(n14697), .Z(n14695) );
  XOR U14540 ( .A(n14583), .B(n14698), .Z(n14577) );
  IV U14541 ( .A(n14582), .Z(n14698) );
  XNOR U14542 ( .A(n14579), .B(n14659), .Z(n14582) );
  AND U14543 ( .A(n15553), .B(n14041), .Z(n14659) );
  XOR U14544 ( .A(n14699), .B(n14700), .Z(n14579) );
  ANDN U14545 ( .A(n14701), .B(n14702), .Z(n14700) );
  XNOR U14546 ( .A(n14699), .B(n14703), .Z(n14701) );
  XOR U14547 ( .A(n14589), .B(n14704), .Z(n14583) );
  IV U14548 ( .A(n14588), .Z(n14704) );
  XNOR U14549 ( .A(n14585), .B(n14652), .Z(n14588) );
  AND U14550 ( .A(n15896), .B(n13880), .Z(n14652) );
  XOR U14551 ( .A(n14705), .B(n14706), .Z(n14585) );
  ANDN U14552 ( .A(n14707), .B(n14708), .Z(n14706) );
  XNOR U14553 ( .A(n14705), .B(n14709), .Z(n14707) );
  XOR U14554 ( .A(n14595), .B(n14710), .Z(n14589) );
  IV U14555 ( .A(n14594), .Z(n14710) );
  XNOR U14556 ( .A(n14591), .B(n14645), .Z(n14594) );
  AND U14557 ( .A(n16265), .B(n13745), .Z(n14645) );
  XOR U14558 ( .A(n14711), .B(n14712), .Z(n14591) );
  ANDN U14559 ( .A(n14713), .B(n14714), .Z(n14712) );
  XNOR U14560 ( .A(n14711), .B(n14715), .Z(n14713) );
  XOR U14561 ( .A(n14601), .B(n14716), .Z(n14595) );
  IV U14562 ( .A(n14600), .Z(n14716) );
  XNOR U14563 ( .A(n14597), .B(n14638), .Z(n14600) );
  AND U14564 ( .A(n16657), .B(n13636), .Z(n14638) );
  XOR U14565 ( .A(n14717), .B(n14718), .Z(n14597) );
  ANDN U14566 ( .A(n14719), .B(n14720), .Z(n14718) );
  XNOR U14567 ( .A(n14717), .B(n14721), .Z(n14719) );
  XOR U14568 ( .A(n14607), .B(n14722), .Z(n14601) );
  IV U14569 ( .A(n14606), .Z(n14722) );
  XNOR U14570 ( .A(n14603), .B(n14631), .Z(n14606) );
  AND U14571 ( .A(n17567), .B(n13553), .Z(n14631) );
  XOR U14572 ( .A(n14723), .B(n14724), .Z(n14603) );
  ANDN U14573 ( .A(n14725), .B(n14726), .Z(n14724) );
  XNOR U14574 ( .A(n14723), .B(n14727), .Z(n14725) );
  XOR U14575 ( .A(n14613), .B(n14728), .Z(n14607) );
  IV U14576 ( .A(n14612), .Z(n14728) );
  XNOR U14577 ( .A(n14609), .B(n14624), .Z(n14612) );
  AND U14578 ( .A(n17688), .B(n13496), .Z(n14624) );
  XOR U14579 ( .A(n14729), .B(n14730), .Z(n14609) );
  ANDN U14580 ( .A(n14731), .B(n14732), .Z(n14730) );
  XNOR U14581 ( .A(n14729), .B(n14733), .Z(n14731) );
  XOR U14582 ( .A(n14618), .B(n14734), .Z(n14613) );
  IV U14583 ( .A(n14617), .Z(n14734) );
  XNOR U14584 ( .A(n14614), .B(n14622), .Z(n14617) );
  AND U14585 ( .A(n13470), .B(n17814), .Z(n14622) );
  XOR U14586 ( .A(n14735), .B(n14736), .Z(n14614) );
  ANDN U14587 ( .A(n14737), .B(n14738), .Z(n14736) );
  XNOR U14588 ( .A(n14735), .B(n14739), .Z(n14737) );
  XNOR U14589 ( .A(n14740), .B(n14741), .Z(n14618) );
  ANDN U14590 ( .A(n14742), .B(n14743), .Z(n14741) );
  XNOR U14591 ( .A(n14740), .B(n14744), .Z(n14742) );
  XOR U14592 ( .A(n14745), .B(n14746), .Z(n14619) );
  ANDN U14593 ( .A(n14747), .B(n6544), .Z(n14746) );
  XNOR U14594 ( .A(n14745), .B(n14748), .Z(n6544) );
  XNOR U14595 ( .A(n14745), .B(n6542), .Z(n14747) );
  XOR U14596 ( .A(n14629), .B(n14749), .Z(n6542) );
  IV U14597 ( .A(n14628), .Z(n14749) );
  XNOR U14598 ( .A(n14625), .B(n14750), .Z(n14628) );
  XOR U14599 ( .A(n14751), .B(n14752), .Z(n14625) );
  ANDN U14600 ( .A(n14753), .B(n14754), .Z(n14752) );
  XNOR U14601 ( .A(n14751), .B(n14755), .Z(n14753) );
  XOR U14602 ( .A(n14636), .B(n14756), .Z(n14629) );
  IV U14603 ( .A(n14635), .Z(n14756) );
  XNOR U14604 ( .A(n14632), .B(n14757), .Z(n14635) );
  XOR U14605 ( .A(n14758), .B(n14759), .Z(n14632) );
  ANDN U14606 ( .A(n14760), .B(n14761), .Z(n14759) );
  XNOR U14607 ( .A(n14758), .B(n14762), .Z(n14760) );
  XOR U14608 ( .A(n14643), .B(n14763), .Z(n14636) );
  IV U14609 ( .A(n14642), .Z(n14763) );
  XNOR U14610 ( .A(n14639), .B(n14764), .Z(n14642) );
  XOR U14611 ( .A(n14765), .B(n14766), .Z(n14639) );
  ANDN U14612 ( .A(n14767), .B(n14768), .Z(n14766) );
  XNOR U14613 ( .A(n14765), .B(n14769), .Z(n14767) );
  XOR U14614 ( .A(n14650), .B(n14770), .Z(n14643) );
  IV U14615 ( .A(n14649), .Z(n14770) );
  XNOR U14616 ( .A(n14646), .B(n14771), .Z(n14649) );
  XOR U14617 ( .A(n14772), .B(n14773), .Z(n14646) );
  ANDN U14618 ( .A(n14774), .B(n14775), .Z(n14773) );
  XNOR U14619 ( .A(n14772), .B(n14776), .Z(n14774) );
  XOR U14620 ( .A(n14657), .B(n14777), .Z(n14650) );
  IV U14621 ( .A(n14656), .Z(n14777) );
  XNOR U14622 ( .A(n14653), .B(n14778), .Z(n14656) );
  XOR U14623 ( .A(n14779), .B(n14780), .Z(n14653) );
  ANDN U14624 ( .A(n14781), .B(n14782), .Z(n14780) );
  XNOR U14625 ( .A(n14779), .B(n14783), .Z(n14781) );
  XOR U14626 ( .A(n14664), .B(n14784), .Z(n14657) );
  IV U14627 ( .A(n14663), .Z(n14784) );
  XNOR U14628 ( .A(n14660), .B(n14785), .Z(n14663) );
  XOR U14629 ( .A(n14786), .B(n14787), .Z(n14660) );
  ANDN U14630 ( .A(n14788), .B(n14789), .Z(n14787) );
  XNOR U14631 ( .A(n14786), .B(n14790), .Z(n14788) );
  XOR U14632 ( .A(n14671), .B(n14791), .Z(n14664) );
  IV U14633 ( .A(n14670), .Z(n14791) );
  XNOR U14634 ( .A(n14667), .B(n14792), .Z(n14670) );
  XOR U14635 ( .A(n14793), .B(n14794), .Z(n14667) );
  ANDN U14636 ( .A(n14795), .B(n14796), .Z(n14794) );
  XNOR U14637 ( .A(n14793), .B(n14797), .Z(n14795) );
  XOR U14638 ( .A(n14678), .B(n14798), .Z(n14671) );
  IV U14639 ( .A(n14677), .Z(n14798) );
  XNOR U14640 ( .A(n14674), .B(n14799), .Z(n14677) );
  XOR U14641 ( .A(n14800), .B(n14801), .Z(n14674) );
  ANDN U14642 ( .A(n14802), .B(n14803), .Z(n14801) );
  XNOR U14643 ( .A(n14800), .B(n14804), .Z(n14802) );
  XOR U14644 ( .A(n14685), .B(n14805), .Z(n14678) );
  IV U14645 ( .A(n14684), .Z(n14805) );
  XNOR U14646 ( .A(n14681), .B(n14806), .Z(n14684) );
  XOR U14647 ( .A(n14807), .B(n14808), .Z(n14681) );
  ANDN U14648 ( .A(n14809), .B(n14810), .Z(n14808) );
  XNOR U14649 ( .A(n14807), .B(n14811), .Z(n14809) );
  XOR U14650 ( .A(n14691), .B(n14812), .Z(n14685) );
  IV U14651 ( .A(n14690), .Z(n14812) );
  XNOR U14652 ( .A(n14687), .B(n14806), .Z(n14690) );
  AND U14653 ( .A(n14945), .B(n14680), .Z(n14806) );
  XOR U14654 ( .A(n14813), .B(n14814), .Z(n14687) );
  ANDN U14655 ( .A(n14815), .B(n14816), .Z(n14814) );
  XNOR U14656 ( .A(n14813), .B(n14817), .Z(n14815) );
  XOR U14657 ( .A(n14697), .B(n14818), .Z(n14691) );
  IV U14658 ( .A(n14696), .Z(n14818) );
  XNOR U14659 ( .A(n14693), .B(n14799), .Z(n14696) );
  AND U14660 ( .A(n15236), .B(n14441), .Z(n14799) );
  XOR U14661 ( .A(n14819), .B(n14820), .Z(n14693) );
  ANDN U14662 ( .A(n14821), .B(n14822), .Z(n14820) );
  XNOR U14663 ( .A(n14819), .B(n14823), .Z(n14821) );
  XOR U14664 ( .A(n14703), .B(n14824), .Z(n14697) );
  IV U14665 ( .A(n14702), .Z(n14824) );
  XNOR U14666 ( .A(n14699), .B(n14792), .Z(n14702) );
  AND U14667 ( .A(n15553), .B(n14228), .Z(n14792) );
  XOR U14668 ( .A(n14825), .B(n14826), .Z(n14699) );
  ANDN U14669 ( .A(n14827), .B(n14828), .Z(n14826) );
  XNOR U14670 ( .A(n14825), .B(n14829), .Z(n14827) );
  XOR U14671 ( .A(n14709), .B(n14830), .Z(n14703) );
  IV U14672 ( .A(n14708), .Z(n14830) );
  XNOR U14673 ( .A(n14705), .B(n14785), .Z(n14708) );
  AND U14674 ( .A(n15896), .B(n14041), .Z(n14785) );
  XOR U14675 ( .A(n14831), .B(n14832), .Z(n14705) );
  ANDN U14676 ( .A(n14833), .B(n14834), .Z(n14832) );
  XNOR U14677 ( .A(n14831), .B(n14835), .Z(n14833) );
  XOR U14678 ( .A(n14715), .B(n14836), .Z(n14709) );
  IV U14679 ( .A(n14714), .Z(n14836) );
  XNOR U14680 ( .A(n14711), .B(n14778), .Z(n14714) );
  AND U14681 ( .A(n16265), .B(n13880), .Z(n14778) );
  XOR U14682 ( .A(n14837), .B(n14838), .Z(n14711) );
  ANDN U14683 ( .A(n14839), .B(n14840), .Z(n14838) );
  XNOR U14684 ( .A(n14837), .B(n14841), .Z(n14839) );
  XOR U14685 ( .A(n14721), .B(n14842), .Z(n14715) );
  IV U14686 ( .A(n14720), .Z(n14842) );
  XNOR U14687 ( .A(n14717), .B(n14771), .Z(n14720) );
  AND U14688 ( .A(n16657), .B(n13745), .Z(n14771) );
  XOR U14689 ( .A(n14843), .B(n14844), .Z(n14717) );
  ANDN U14690 ( .A(n14845), .B(n14846), .Z(n14844) );
  XNOR U14691 ( .A(n14843), .B(n14847), .Z(n14845) );
  XOR U14692 ( .A(n14727), .B(n14848), .Z(n14721) );
  IV U14693 ( .A(n14726), .Z(n14848) );
  XNOR U14694 ( .A(n14723), .B(n14764), .Z(n14726) );
  AND U14695 ( .A(n17567), .B(n13636), .Z(n14764) );
  XOR U14696 ( .A(n14849), .B(n14850), .Z(n14723) );
  ANDN U14697 ( .A(n14851), .B(n14852), .Z(n14850) );
  XNOR U14698 ( .A(n14849), .B(n14853), .Z(n14851) );
  XOR U14699 ( .A(n14733), .B(n14854), .Z(n14727) );
  IV U14700 ( .A(n14732), .Z(n14854) );
  XNOR U14701 ( .A(n14729), .B(n14757), .Z(n14732) );
  AND U14702 ( .A(n17688), .B(n13553), .Z(n14757) );
  XOR U14703 ( .A(n14855), .B(n14856), .Z(n14729) );
  ANDN U14704 ( .A(n14857), .B(n14858), .Z(n14856) );
  XNOR U14705 ( .A(n14855), .B(n14859), .Z(n14857) );
  XOR U14706 ( .A(n14739), .B(n14860), .Z(n14733) );
  IV U14707 ( .A(n14738), .Z(n14860) );
  XNOR U14708 ( .A(n14735), .B(n14750), .Z(n14738) );
  AND U14709 ( .A(n17814), .B(n13496), .Z(n14750) );
  XOR U14710 ( .A(n14861), .B(n14862), .Z(n14735) );
  ANDN U14711 ( .A(n14863), .B(n14864), .Z(n14862) );
  XNOR U14712 ( .A(n14861), .B(n14865), .Z(n14863) );
  XOR U14713 ( .A(n14744), .B(n14866), .Z(n14739) );
  IV U14714 ( .A(n14743), .Z(n14866) );
  XNOR U14715 ( .A(n14740), .B(n14748), .Z(n14743) );
  AND U14716 ( .A(n13470), .B(n17945), .Z(n14748) );
  XOR U14717 ( .A(n14867), .B(n14868), .Z(n14740) );
  ANDN U14718 ( .A(n14869), .B(n14870), .Z(n14868) );
  XNOR U14719 ( .A(n14867), .B(n14871), .Z(n14869) );
  XNOR U14720 ( .A(n14872), .B(n14873), .Z(n14744) );
  ANDN U14721 ( .A(n14874), .B(n14875), .Z(n14873) );
  XNOR U14722 ( .A(n14872), .B(n14876), .Z(n14874) );
  XOR U14723 ( .A(n14877), .B(n14878), .Z(n14745) );
  ANDN U14724 ( .A(n14879), .B(n6828), .Z(n14878) );
  XNOR U14725 ( .A(n14877), .B(n14880), .Z(n6828) );
  XNOR U14726 ( .A(n14877), .B(n6826), .Z(n14879) );
  XOR U14727 ( .A(n14755), .B(n14881), .Z(n6826) );
  IV U14728 ( .A(n14754), .Z(n14881) );
  XNOR U14729 ( .A(n14751), .B(n14882), .Z(n14754) );
  XOR U14730 ( .A(n14883), .B(n14884), .Z(n14751) );
  ANDN U14731 ( .A(n14885), .B(n14886), .Z(n14884) );
  XNOR U14732 ( .A(n14883), .B(n14887), .Z(n14885) );
  XOR U14733 ( .A(n14762), .B(n14888), .Z(n14755) );
  IV U14734 ( .A(n14761), .Z(n14888) );
  XNOR U14735 ( .A(n14758), .B(n14889), .Z(n14761) );
  XOR U14736 ( .A(n14890), .B(n14891), .Z(n14758) );
  ANDN U14737 ( .A(n14892), .B(n14893), .Z(n14891) );
  XNOR U14738 ( .A(n14890), .B(n14894), .Z(n14892) );
  XOR U14739 ( .A(n14769), .B(n14895), .Z(n14762) );
  IV U14740 ( .A(n14768), .Z(n14895) );
  XNOR U14741 ( .A(n14765), .B(n14896), .Z(n14768) );
  XOR U14742 ( .A(n14897), .B(n14898), .Z(n14765) );
  ANDN U14743 ( .A(n14899), .B(n14900), .Z(n14898) );
  XNOR U14744 ( .A(n14897), .B(n14901), .Z(n14899) );
  XOR U14745 ( .A(n14776), .B(n14902), .Z(n14769) );
  IV U14746 ( .A(n14775), .Z(n14902) );
  XNOR U14747 ( .A(n14772), .B(n14903), .Z(n14775) );
  XOR U14748 ( .A(n14904), .B(n14905), .Z(n14772) );
  ANDN U14749 ( .A(n14906), .B(n14907), .Z(n14905) );
  XNOR U14750 ( .A(n14904), .B(n14908), .Z(n14906) );
  XOR U14751 ( .A(n14783), .B(n14909), .Z(n14776) );
  IV U14752 ( .A(n14782), .Z(n14909) );
  XNOR U14753 ( .A(n14779), .B(n14910), .Z(n14782) );
  XOR U14754 ( .A(n14911), .B(n14912), .Z(n14779) );
  ANDN U14755 ( .A(n14913), .B(n14914), .Z(n14912) );
  XNOR U14756 ( .A(n14911), .B(n14915), .Z(n14913) );
  XOR U14757 ( .A(n14790), .B(n14916), .Z(n14783) );
  IV U14758 ( .A(n14789), .Z(n14916) );
  XNOR U14759 ( .A(n14786), .B(n14917), .Z(n14789) );
  XOR U14760 ( .A(n14918), .B(n14919), .Z(n14786) );
  ANDN U14761 ( .A(n14920), .B(n14921), .Z(n14919) );
  XNOR U14762 ( .A(n14918), .B(n14922), .Z(n14920) );
  XOR U14763 ( .A(n14797), .B(n14923), .Z(n14790) );
  IV U14764 ( .A(n14796), .Z(n14923) );
  XNOR U14765 ( .A(n14793), .B(n14924), .Z(n14796) );
  XOR U14766 ( .A(n14925), .B(n14926), .Z(n14793) );
  ANDN U14767 ( .A(n14927), .B(n14928), .Z(n14926) );
  XNOR U14768 ( .A(n14925), .B(n14929), .Z(n14927) );
  XOR U14769 ( .A(n14804), .B(n14930), .Z(n14797) );
  IV U14770 ( .A(n14803), .Z(n14930) );
  XNOR U14771 ( .A(n14800), .B(n14931), .Z(n14803) );
  XOR U14772 ( .A(n14932), .B(n14933), .Z(n14800) );
  ANDN U14773 ( .A(n14934), .B(n14935), .Z(n14933) );
  XNOR U14774 ( .A(n14932), .B(n14936), .Z(n14934) );
  XOR U14775 ( .A(n14811), .B(n14937), .Z(n14804) );
  IV U14776 ( .A(n14810), .Z(n14937) );
  XNOR U14777 ( .A(n14807), .B(n14938), .Z(n14810) );
  XOR U14778 ( .A(n14939), .B(n14940), .Z(n14807) );
  ANDN U14779 ( .A(n14941), .B(n14942), .Z(n14940) );
  XNOR U14780 ( .A(n14939), .B(n14943), .Z(n14941) );
  XOR U14781 ( .A(n14817), .B(n14944), .Z(n14811) );
  IV U14782 ( .A(n14816), .Z(n14944) );
  XNOR U14783 ( .A(n14813), .B(n14945), .Z(n14816) );
  XOR U14784 ( .A(n14946), .B(n14947), .Z(n14813) );
  ANDN U14785 ( .A(n14948), .B(n14949), .Z(n14947) );
  XNOR U14786 ( .A(n14946), .B(n14950), .Z(n14948) );
  XOR U14787 ( .A(n14823), .B(n14951), .Z(n14817) );
  IV U14788 ( .A(n14822), .Z(n14951) );
  XNOR U14789 ( .A(n14819), .B(n14938), .Z(n14822) );
  AND U14790 ( .A(n15236), .B(n14680), .Z(n14938) );
  XOR U14791 ( .A(n14952), .B(n14953), .Z(n14819) );
  ANDN U14792 ( .A(n14954), .B(n14955), .Z(n14953) );
  XNOR U14793 ( .A(n14952), .B(n14956), .Z(n14954) );
  XOR U14794 ( .A(n14829), .B(n14957), .Z(n14823) );
  IV U14795 ( .A(n14828), .Z(n14957) );
  XNOR U14796 ( .A(n14825), .B(n14931), .Z(n14828) );
  AND U14797 ( .A(n15553), .B(n14441), .Z(n14931) );
  XOR U14798 ( .A(n14958), .B(n14959), .Z(n14825) );
  ANDN U14799 ( .A(n14960), .B(n14961), .Z(n14959) );
  XNOR U14800 ( .A(n14958), .B(n14962), .Z(n14960) );
  XOR U14801 ( .A(n14835), .B(n14963), .Z(n14829) );
  IV U14802 ( .A(n14834), .Z(n14963) );
  XNOR U14803 ( .A(n14831), .B(n14924), .Z(n14834) );
  AND U14804 ( .A(n15896), .B(n14228), .Z(n14924) );
  XOR U14805 ( .A(n14964), .B(n14965), .Z(n14831) );
  ANDN U14806 ( .A(n14966), .B(n14967), .Z(n14965) );
  XNOR U14807 ( .A(n14964), .B(n14968), .Z(n14966) );
  XOR U14808 ( .A(n14841), .B(n14969), .Z(n14835) );
  IV U14809 ( .A(n14840), .Z(n14969) );
  XNOR U14810 ( .A(n14837), .B(n14917), .Z(n14840) );
  AND U14811 ( .A(n16265), .B(n14041), .Z(n14917) );
  XOR U14812 ( .A(n14970), .B(n14971), .Z(n14837) );
  ANDN U14813 ( .A(n14972), .B(n14973), .Z(n14971) );
  XNOR U14814 ( .A(n14970), .B(n14974), .Z(n14972) );
  XOR U14815 ( .A(n14847), .B(n14975), .Z(n14841) );
  IV U14816 ( .A(n14846), .Z(n14975) );
  XNOR U14817 ( .A(n14843), .B(n14910), .Z(n14846) );
  AND U14818 ( .A(n16657), .B(n13880), .Z(n14910) );
  XOR U14819 ( .A(n14976), .B(n14977), .Z(n14843) );
  ANDN U14820 ( .A(n14978), .B(n14979), .Z(n14977) );
  XNOR U14821 ( .A(n14976), .B(n14980), .Z(n14978) );
  XOR U14822 ( .A(n14853), .B(n14981), .Z(n14847) );
  IV U14823 ( .A(n14852), .Z(n14981) );
  XNOR U14824 ( .A(n14849), .B(n14903), .Z(n14852) );
  AND U14825 ( .A(n17567), .B(n13745), .Z(n14903) );
  XOR U14826 ( .A(n14982), .B(n14983), .Z(n14849) );
  ANDN U14827 ( .A(n14984), .B(n14985), .Z(n14983) );
  XNOR U14828 ( .A(n14982), .B(n14986), .Z(n14984) );
  XOR U14829 ( .A(n14859), .B(n14987), .Z(n14853) );
  IV U14830 ( .A(n14858), .Z(n14987) );
  XNOR U14831 ( .A(n14855), .B(n14896), .Z(n14858) );
  AND U14832 ( .A(n17688), .B(n13636), .Z(n14896) );
  XOR U14833 ( .A(n14988), .B(n14989), .Z(n14855) );
  ANDN U14834 ( .A(n14990), .B(n14991), .Z(n14989) );
  XNOR U14835 ( .A(n14988), .B(n14992), .Z(n14990) );
  XOR U14836 ( .A(n14865), .B(n14993), .Z(n14859) );
  IV U14837 ( .A(n14864), .Z(n14993) );
  XNOR U14838 ( .A(n14861), .B(n14889), .Z(n14864) );
  AND U14839 ( .A(n17814), .B(n13553), .Z(n14889) );
  XOR U14840 ( .A(n14994), .B(n14995), .Z(n14861) );
  ANDN U14841 ( .A(n14996), .B(n14997), .Z(n14995) );
  XNOR U14842 ( .A(n14994), .B(n14998), .Z(n14996) );
  XOR U14843 ( .A(n14871), .B(n14999), .Z(n14865) );
  IV U14844 ( .A(n14870), .Z(n14999) );
  XNOR U14845 ( .A(n14867), .B(n14882), .Z(n14870) );
  AND U14846 ( .A(n17945), .B(n13496), .Z(n14882) );
  XOR U14847 ( .A(n15000), .B(n15001), .Z(n14867) );
  ANDN U14848 ( .A(n15002), .B(n15003), .Z(n15001) );
  XNOR U14849 ( .A(n15000), .B(n15004), .Z(n15002) );
  XOR U14850 ( .A(n14876), .B(n15005), .Z(n14871) );
  IV U14851 ( .A(n14875), .Z(n15005) );
  XNOR U14852 ( .A(n14872), .B(n14880), .Z(n14875) );
  AND U14853 ( .A(n13470), .B(n18081), .Z(n14880) );
  XOR U14854 ( .A(n15006), .B(n15007), .Z(n14872) );
  ANDN U14855 ( .A(n15008), .B(n15009), .Z(n15007) );
  XNOR U14856 ( .A(n15006), .B(n15010), .Z(n15008) );
  XNOR U14857 ( .A(n15011), .B(n15012), .Z(n14876) );
  ANDN U14858 ( .A(n15013), .B(n15014), .Z(n15012) );
  XNOR U14859 ( .A(n15011), .B(n15015), .Z(n15013) );
  XOR U14860 ( .A(n15016), .B(n15017), .Z(n14877) );
  ANDN U14861 ( .A(n15018), .B(n7104), .Z(n15017) );
  XNOR U14862 ( .A(n15016), .B(n15019), .Z(n7104) );
  XNOR U14863 ( .A(n15016), .B(n7102), .Z(n15018) );
  XOR U14864 ( .A(n14887), .B(n15020), .Z(n7102) );
  IV U14865 ( .A(n14886), .Z(n15020) );
  XNOR U14866 ( .A(n14883), .B(n15021), .Z(n14886) );
  XOR U14867 ( .A(n15022), .B(n15023), .Z(n14883) );
  ANDN U14868 ( .A(n15024), .B(n15025), .Z(n15023) );
  XNOR U14869 ( .A(n15022), .B(n15026), .Z(n15024) );
  XOR U14870 ( .A(n14894), .B(n15027), .Z(n14887) );
  IV U14871 ( .A(n14893), .Z(n15027) );
  XNOR U14872 ( .A(n14890), .B(n15028), .Z(n14893) );
  XOR U14873 ( .A(n15029), .B(n15030), .Z(n14890) );
  ANDN U14874 ( .A(n15031), .B(n15032), .Z(n15030) );
  XNOR U14875 ( .A(n15029), .B(n15033), .Z(n15031) );
  XOR U14876 ( .A(n14901), .B(n15034), .Z(n14894) );
  IV U14877 ( .A(n14900), .Z(n15034) );
  XNOR U14878 ( .A(n14897), .B(n15035), .Z(n14900) );
  XOR U14879 ( .A(n15036), .B(n15037), .Z(n14897) );
  ANDN U14880 ( .A(n15038), .B(n15039), .Z(n15037) );
  XNOR U14881 ( .A(n15036), .B(n15040), .Z(n15038) );
  XOR U14882 ( .A(n14908), .B(n15041), .Z(n14901) );
  IV U14883 ( .A(n14907), .Z(n15041) );
  XNOR U14884 ( .A(n14904), .B(n15042), .Z(n14907) );
  XOR U14885 ( .A(n15043), .B(n15044), .Z(n14904) );
  ANDN U14886 ( .A(n15045), .B(n15046), .Z(n15044) );
  XNOR U14887 ( .A(n15043), .B(n15047), .Z(n15045) );
  XOR U14888 ( .A(n14915), .B(n15048), .Z(n14908) );
  IV U14889 ( .A(n14914), .Z(n15048) );
  XNOR U14890 ( .A(n14911), .B(n15049), .Z(n14914) );
  XOR U14891 ( .A(n15050), .B(n15051), .Z(n14911) );
  ANDN U14892 ( .A(n15052), .B(n15053), .Z(n15051) );
  XNOR U14893 ( .A(n15050), .B(n15054), .Z(n15052) );
  XOR U14894 ( .A(n14922), .B(n15055), .Z(n14915) );
  IV U14895 ( .A(n14921), .Z(n15055) );
  XNOR U14896 ( .A(n14918), .B(n15056), .Z(n14921) );
  XOR U14897 ( .A(n15057), .B(n15058), .Z(n14918) );
  ANDN U14898 ( .A(n15059), .B(n15060), .Z(n15058) );
  XNOR U14899 ( .A(n15057), .B(n15061), .Z(n15059) );
  XOR U14900 ( .A(n14929), .B(n15062), .Z(n14922) );
  IV U14901 ( .A(n14928), .Z(n15062) );
  XNOR U14902 ( .A(n14925), .B(n15063), .Z(n14928) );
  XOR U14903 ( .A(n15064), .B(n15065), .Z(n14925) );
  ANDN U14904 ( .A(n15066), .B(n15067), .Z(n15065) );
  XNOR U14905 ( .A(n15064), .B(n15068), .Z(n15066) );
  XOR U14906 ( .A(n14936), .B(n15069), .Z(n14929) );
  IV U14907 ( .A(n14935), .Z(n15069) );
  XNOR U14908 ( .A(n14932), .B(n15070), .Z(n14935) );
  XOR U14909 ( .A(n15071), .B(n15072), .Z(n14932) );
  ANDN U14910 ( .A(n15073), .B(n15074), .Z(n15072) );
  XNOR U14911 ( .A(n15071), .B(n15075), .Z(n15073) );
  XOR U14912 ( .A(n14943), .B(n15076), .Z(n14936) );
  IV U14913 ( .A(n14942), .Z(n15076) );
  XNOR U14914 ( .A(n14939), .B(n15077), .Z(n14942) );
  XOR U14915 ( .A(n15078), .B(n15079), .Z(n14939) );
  ANDN U14916 ( .A(n15080), .B(n15081), .Z(n15079) );
  XNOR U14917 ( .A(n15078), .B(n15082), .Z(n15080) );
  XOR U14918 ( .A(n14950), .B(n15083), .Z(n14943) );
  IV U14919 ( .A(n14949), .Z(n15083) );
  XNOR U14920 ( .A(n14946), .B(n15084), .Z(n14949) );
  XOR U14921 ( .A(n15085), .B(n15086), .Z(n14946) );
  ANDN U14922 ( .A(n15087), .B(n15088), .Z(n15086) );
  XNOR U14923 ( .A(n15085), .B(n15089), .Z(n15087) );
  XOR U14924 ( .A(n14956), .B(n15090), .Z(n14950) );
  IV U14925 ( .A(n14955), .Z(n15090) );
  XNOR U14926 ( .A(n14952), .B(n15084), .Z(n14955) );
  AND U14927 ( .A(n15236), .B(n14945), .Z(n15084) );
  XOR U14928 ( .A(n15091), .B(n15092), .Z(n14952) );
  ANDN U14929 ( .A(n15093), .B(n15094), .Z(n15092) );
  XNOR U14930 ( .A(n15091), .B(n15095), .Z(n15093) );
  XOR U14931 ( .A(n14962), .B(n15096), .Z(n14956) );
  IV U14932 ( .A(n14961), .Z(n15096) );
  XNOR U14933 ( .A(n14958), .B(n15077), .Z(n14961) );
  AND U14934 ( .A(n15553), .B(n14680), .Z(n15077) );
  XOR U14935 ( .A(n15097), .B(n15098), .Z(n14958) );
  ANDN U14936 ( .A(n15099), .B(n15100), .Z(n15098) );
  XNOR U14937 ( .A(n15097), .B(n15101), .Z(n15099) );
  XOR U14938 ( .A(n14968), .B(n15102), .Z(n14962) );
  IV U14939 ( .A(n14967), .Z(n15102) );
  XNOR U14940 ( .A(n14964), .B(n15070), .Z(n14967) );
  AND U14941 ( .A(n15896), .B(n14441), .Z(n15070) );
  XOR U14942 ( .A(n15103), .B(n15104), .Z(n14964) );
  ANDN U14943 ( .A(n15105), .B(n15106), .Z(n15104) );
  XNOR U14944 ( .A(n15103), .B(n15107), .Z(n15105) );
  XOR U14945 ( .A(n14974), .B(n15108), .Z(n14968) );
  IV U14946 ( .A(n14973), .Z(n15108) );
  XNOR U14947 ( .A(n14970), .B(n15063), .Z(n14973) );
  AND U14948 ( .A(n16265), .B(n14228), .Z(n15063) );
  XOR U14949 ( .A(n15109), .B(n15110), .Z(n14970) );
  ANDN U14950 ( .A(n15111), .B(n15112), .Z(n15110) );
  XNOR U14951 ( .A(n15109), .B(n15113), .Z(n15111) );
  XOR U14952 ( .A(n14980), .B(n15114), .Z(n14974) );
  IV U14953 ( .A(n14979), .Z(n15114) );
  XNOR U14954 ( .A(n14976), .B(n15056), .Z(n14979) );
  AND U14955 ( .A(n16657), .B(n14041), .Z(n15056) );
  XOR U14956 ( .A(n15115), .B(n15116), .Z(n14976) );
  ANDN U14957 ( .A(n15117), .B(n15118), .Z(n15116) );
  XNOR U14958 ( .A(n15115), .B(n15119), .Z(n15117) );
  XOR U14959 ( .A(n14986), .B(n15120), .Z(n14980) );
  IV U14960 ( .A(n14985), .Z(n15120) );
  XNOR U14961 ( .A(n14982), .B(n15049), .Z(n14985) );
  AND U14962 ( .A(n17567), .B(n13880), .Z(n15049) );
  XOR U14963 ( .A(n15121), .B(n15122), .Z(n14982) );
  ANDN U14964 ( .A(n15123), .B(n15124), .Z(n15122) );
  XNOR U14965 ( .A(n15121), .B(n15125), .Z(n15123) );
  XOR U14966 ( .A(n14992), .B(n15126), .Z(n14986) );
  IV U14967 ( .A(n14991), .Z(n15126) );
  XNOR U14968 ( .A(n14988), .B(n15042), .Z(n14991) );
  AND U14969 ( .A(n17688), .B(n13745), .Z(n15042) );
  XOR U14970 ( .A(n15127), .B(n15128), .Z(n14988) );
  ANDN U14971 ( .A(n15129), .B(n15130), .Z(n15128) );
  XNOR U14972 ( .A(n15127), .B(n15131), .Z(n15129) );
  XOR U14973 ( .A(n14998), .B(n15132), .Z(n14992) );
  IV U14974 ( .A(n14997), .Z(n15132) );
  XNOR U14975 ( .A(n14994), .B(n15035), .Z(n14997) );
  AND U14976 ( .A(n17814), .B(n13636), .Z(n15035) );
  XOR U14977 ( .A(n15133), .B(n15134), .Z(n14994) );
  ANDN U14978 ( .A(n15135), .B(n15136), .Z(n15134) );
  XNOR U14979 ( .A(n15133), .B(n15137), .Z(n15135) );
  XOR U14980 ( .A(n15004), .B(n15138), .Z(n14998) );
  IV U14981 ( .A(n15003), .Z(n15138) );
  XNOR U14982 ( .A(n15000), .B(n15028), .Z(n15003) );
  AND U14983 ( .A(n17945), .B(n13553), .Z(n15028) );
  XOR U14984 ( .A(n15139), .B(n15140), .Z(n15000) );
  ANDN U14985 ( .A(n15141), .B(n15142), .Z(n15140) );
  XNOR U14986 ( .A(n15139), .B(n15143), .Z(n15141) );
  XOR U14987 ( .A(n15010), .B(n15144), .Z(n15004) );
  IV U14988 ( .A(n15009), .Z(n15144) );
  XNOR U14989 ( .A(n15006), .B(n15021), .Z(n15009) );
  AND U14990 ( .A(n18081), .B(n13496), .Z(n15021) );
  XOR U14991 ( .A(n15145), .B(n15146), .Z(n15006) );
  ANDN U14992 ( .A(n15147), .B(n15148), .Z(n15146) );
  XNOR U14993 ( .A(n15145), .B(n15149), .Z(n15147) );
  XOR U14994 ( .A(n15015), .B(n15150), .Z(n15010) );
  IV U14995 ( .A(n15014), .Z(n15150) );
  XNOR U14996 ( .A(n15011), .B(n15019), .Z(n15014) );
  AND U14997 ( .A(n13470), .B(n18222), .Z(n15019) );
  XOR U14998 ( .A(n15151), .B(n15152), .Z(n15011) );
  ANDN U14999 ( .A(n15153), .B(n15154), .Z(n15152) );
  XNOR U15000 ( .A(n15151), .B(n15155), .Z(n15153) );
  XNOR U15001 ( .A(n15156), .B(n15157), .Z(n15015) );
  ANDN U15002 ( .A(n15158), .B(n15159), .Z(n15157) );
  XNOR U15003 ( .A(n15156), .B(n15160), .Z(n15158) );
  XOR U15004 ( .A(n15161), .B(n15162), .Z(n15016) );
  ANDN U15005 ( .A(n15163), .B(n7376), .Z(n15162) );
  XNOR U15006 ( .A(n15161), .B(n15164), .Z(n7376) );
  XNOR U15007 ( .A(n15161), .B(n7374), .Z(n15163) );
  XOR U15008 ( .A(n15026), .B(n15165), .Z(n7374) );
  IV U15009 ( .A(n15025), .Z(n15165) );
  XNOR U15010 ( .A(n15022), .B(n15166), .Z(n15025) );
  XOR U15011 ( .A(n15167), .B(n15168), .Z(n15022) );
  ANDN U15012 ( .A(n15169), .B(n15170), .Z(n15168) );
  XNOR U15013 ( .A(n15167), .B(n15171), .Z(n15169) );
  XOR U15014 ( .A(n15033), .B(n15172), .Z(n15026) );
  IV U15015 ( .A(n15032), .Z(n15172) );
  XNOR U15016 ( .A(n15029), .B(n15173), .Z(n15032) );
  XOR U15017 ( .A(n15174), .B(n15175), .Z(n15029) );
  ANDN U15018 ( .A(n15176), .B(n15177), .Z(n15175) );
  XNOR U15019 ( .A(n15174), .B(n15178), .Z(n15176) );
  XOR U15020 ( .A(n15040), .B(n15179), .Z(n15033) );
  IV U15021 ( .A(n15039), .Z(n15179) );
  XNOR U15022 ( .A(n15036), .B(n15180), .Z(n15039) );
  XOR U15023 ( .A(n15181), .B(n15182), .Z(n15036) );
  ANDN U15024 ( .A(n15183), .B(n15184), .Z(n15182) );
  XNOR U15025 ( .A(n15181), .B(n15185), .Z(n15183) );
  XOR U15026 ( .A(n15047), .B(n15186), .Z(n15040) );
  IV U15027 ( .A(n15046), .Z(n15186) );
  XNOR U15028 ( .A(n15043), .B(n15187), .Z(n15046) );
  XOR U15029 ( .A(n15188), .B(n15189), .Z(n15043) );
  ANDN U15030 ( .A(n15190), .B(n15191), .Z(n15189) );
  XNOR U15031 ( .A(n15188), .B(n15192), .Z(n15190) );
  XOR U15032 ( .A(n15054), .B(n15193), .Z(n15047) );
  IV U15033 ( .A(n15053), .Z(n15193) );
  XNOR U15034 ( .A(n15050), .B(n15194), .Z(n15053) );
  XOR U15035 ( .A(n15195), .B(n15196), .Z(n15050) );
  ANDN U15036 ( .A(n15197), .B(n15198), .Z(n15196) );
  XNOR U15037 ( .A(n15195), .B(n15199), .Z(n15197) );
  XOR U15038 ( .A(n15061), .B(n15200), .Z(n15054) );
  IV U15039 ( .A(n15060), .Z(n15200) );
  XNOR U15040 ( .A(n15057), .B(n15201), .Z(n15060) );
  XOR U15041 ( .A(n15202), .B(n15203), .Z(n15057) );
  ANDN U15042 ( .A(n15204), .B(n15205), .Z(n15203) );
  XNOR U15043 ( .A(n15202), .B(n15206), .Z(n15204) );
  XOR U15044 ( .A(n15068), .B(n15207), .Z(n15061) );
  IV U15045 ( .A(n15067), .Z(n15207) );
  XNOR U15046 ( .A(n15064), .B(n15208), .Z(n15067) );
  XOR U15047 ( .A(n15209), .B(n15210), .Z(n15064) );
  ANDN U15048 ( .A(n15211), .B(n15212), .Z(n15210) );
  XNOR U15049 ( .A(n15209), .B(n15213), .Z(n15211) );
  XOR U15050 ( .A(n15075), .B(n15214), .Z(n15068) );
  IV U15051 ( .A(n15074), .Z(n15214) );
  XNOR U15052 ( .A(n15071), .B(n15215), .Z(n15074) );
  XOR U15053 ( .A(n15216), .B(n15217), .Z(n15071) );
  ANDN U15054 ( .A(n15218), .B(n15219), .Z(n15217) );
  XNOR U15055 ( .A(n15216), .B(n15220), .Z(n15218) );
  XOR U15056 ( .A(n15082), .B(n15221), .Z(n15075) );
  IV U15057 ( .A(n15081), .Z(n15221) );
  XNOR U15058 ( .A(n15078), .B(n15222), .Z(n15081) );
  XOR U15059 ( .A(n15223), .B(n15224), .Z(n15078) );
  ANDN U15060 ( .A(n15225), .B(n15226), .Z(n15224) );
  XNOR U15061 ( .A(n15223), .B(n15227), .Z(n15225) );
  XOR U15062 ( .A(n15089), .B(n15228), .Z(n15082) );
  IV U15063 ( .A(n15088), .Z(n15228) );
  XNOR U15064 ( .A(n15085), .B(n15229), .Z(n15088) );
  XOR U15065 ( .A(n15230), .B(n15231), .Z(n15085) );
  ANDN U15066 ( .A(n15232), .B(n15233), .Z(n15231) );
  XNOR U15067 ( .A(n15230), .B(n15234), .Z(n15232) );
  XOR U15068 ( .A(n15095), .B(n15235), .Z(n15089) );
  IV U15069 ( .A(n15094), .Z(n15235) );
  XNOR U15070 ( .A(n15091), .B(n15236), .Z(n15094) );
  XOR U15071 ( .A(n15237), .B(n15238), .Z(n15091) );
  ANDN U15072 ( .A(n15239), .B(n15240), .Z(n15238) );
  XNOR U15073 ( .A(n15237), .B(n15241), .Z(n15239) );
  XOR U15074 ( .A(n15101), .B(n15242), .Z(n15095) );
  IV U15075 ( .A(n15100), .Z(n15242) );
  XNOR U15076 ( .A(n15097), .B(n15229), .Z(n15100) );
  AND U15077 ( .A(n15553), .B(n14945), .Z(n15229) );
  XOR U15078 ( .A(n15243), .B(n15244), .Z(n15097) );
  ANDN U15079 ( .A(n15245), .B(n15246), .Z(n15244) );
  XNOR U15080 ( .A(n15243), .B(n15247), .Z(n15245) );
  XOR U15081 ( .A(n15107), .B(n15248), .Z(n15101) );
  IV U15082 ( .A(n15106), .Z(n15248) );
  XNOR U15083 ( .A(n15103), .B(n15222), .Z(n15106) );
  AND U15084 ( .A(n15896), .B(n14680), .Z(n15222) );
  XOR U15085 ( .A(n15249), .B(n15250), .Z(n15103) );
  ANDN U15086 ( .A(n15251), .B(n15252), .Z(n15250) );
  XNOR U15087 ( .A(n15249), .B(n15253), .Z(n15251) );
  XOR U15088 ( .A(n15113), .B(n15254), .Z(n15107) );
  IV U15089 ( .A(n15112), .Z(n15254) );
  XNOR U15090 ( .A(n15109), .B(n15215), .Z(n15112) );
  AND U15091 ( .A(n16265), .B(n14441), .Z(n15215) );
  XOR U15092 ( .A(n15255), .B(n15256), .Z(n15109) );
  ANDN U15093 ( .A(n15257), .B(n15258), .Z(n15256) );
  XNOR U15094 ( .A(n15255), .B(n15259), .Z(n15257) );
  XOR U15095 ( .A(n15119), .B(n15260), .Z(n15113) );
  IV U15096 ( .A(n15118), .Z(n15260) );
  XNOR U15097 ( .A(n15115), .B(n15208), .Z(n15118) );
  AND U15098 ( .A(n16657), .B(n14228), .Z(n15208) );
  XOR U15099 ( .A(n15261), .B(n15262), .Z(n15115) );
  ANDN U15100 ( .A(n15263), .B(n15264), .Z(n15262) );
  XNOR U15101 ( .A(n15261), .B(n15265), .Z(n15263) );
  XOR U15102 ( .A(n15125), .B(n15266), .Z(n15119) );
  IV U15103 ( .A(n15124), .Z(n15266) );
  XNOR U15104 ( .A(n15121), .B(n15201), .Z(n15124) );
  AND U15105 ( .A(n17567), .B(n14041), .Z(n15201) );
  XOR U15106 ( .A(n15267), .B(n15268), .Z(n15121) );
  ANDN U15107 ( .A(n15269), .B(n15270), .Z(n15268) );
  XNOR U15108 ( .A(n15267), .B(n15271), .Z(n15269) );
  XOR U15109 ( .A(n15131), .B(n15272), .Z(n15125) );
  IV U15110 ( .A(n15130), .Z(n15272) );
  XNOR U15111 ( .A(n15127), .B(n15194), .Z(n15130) );
  AND U15112 ( .A(n17688), .B(n13880), .Z(n15194) );
  XOR U15113 ( .A(n15273), .B(n15274), .Z(n15127) );
  ANDN U15114 ( .A(n15275), .B(n15276), .Z(n15274) );
  XNOR U15115 ( .A(n15273), .B(n15277), .Z(n15275) );
  XOR U15116 ( .A(n15137), .B(n15278), .Z(n15131) );
  IV U15117 ( .A(n15136), .Z(n15278) );
  XNOR U15118 ( .A(n15133), .B(n15187), .Z(n15136) );
  AND U15119 ( .A(n17814), .B(n13745), .Z(n15187) );
  XOR U15120 ( .A(n15279), .B(n15280), .Z(n15133) );
  ANDN U15121 ( .A(n15281), .B(n15282), .Z(n15280) );
  XNOR U15122 ( .A(n15279), .B(n15283), .Z(n15281) );
  XOR U15123 ( .A(n15143), .B(n15284), .Z(n15137) );
  IV U15124 ( .A(n15142), .Z(n15284) );
  XNOR U15125 ( .A(n15139), .B(n15180), .Z(n15142) );
  AND U15126 ( .A(n17945), .B(n13636), .Z(n15180) );
  XOR U15127 ( .A(n15285), .B(n15286), .Z(n15139) );
  ANDN U15128 ( .A(n15287), .B(n15288), .Z(n15286) );
  XNOR U15129 ( .A(n15285), .B(n15289), .Z(n15287) );
  XOR U15130 ( .A(n15149), .B(n15290), .Z(n15143) );
  IV U15131 ( .A(n15148), .Z(n15290) );
  XNOR U15132 ( .A(n15145), .B(n15173), .Z(n15148) );
  AND U15133 ( .A(n18081), .B(n13553), .Z(n15173) );
  XOR U15134 ( .A(n15291), .B(n15292), .Z(n15145) );
  ANDN U15135 ( .A(n15293), .B(n15294), .Z(n15292) );
  XNOR U15136 ( .A(n15291), .B(n15295), .Z(n15293) );
  XOR U15137 ( .A(n15155), .B(n15296), .Z(n15149) );
  IV U15138 ( .A(n15154), .Z(n15296) );
  XNOR U15139 ( .A(n15151), .B(n15166), .Z(n15154) );
  AND U15140 ( .A(n18222), .B(n13496), .Z(n15166) );
  XOR U15141 ( .A(n15297), .B(n15298), .Z(n15151) );
  ANDN U15142 ( .A(n15299), .B(n15300), .Z(n15298) );
  XNOR U15143 ( .A(n15297), .B(n15301), .Z(n15299) );
  XOR U15144 ( .A(n15160), .B(n15302), .Z(n15155) );
  IV U15145 ( .A(n15159), .Z(n15302) );
  XNOR U15146 ( .A(n15156), .B(n15164), .Z(n15159) );
  AND U15147 ( .A(n13470), .B(n18368), .Z(n15164) );
  XOR U15148 ( .A(n15303), .B(n15304), .Z(n15156) );
  ANDN U15149 ( .A(n15305), .B(n15306), .Z(n15304) );
  XNOR U15150 ( .A(n15303), .B(n15307), .Z(n15305) );
  XNOR U15151 ( .A(n15308), .B(n15309), .Z(n15160) );
  ANDN U15152 ( .A(n15310), .B(n15311), .Z(n15309) );
  XNOR U15153 ( .A(n15308), .B(n15312), .Z(n15310) );
  XOR U15154 ( .A(n15313), .B(n15314), .Z(n15161) );
  ANDN U15155 ( .A(n15315), .B(n7640), .Z(n15314) );
  XNOR U15156 ( .A(n15313), .B(n15316), .Z(n7640) );
  XNOR U15157 ( .A(n15313), .B(n7638), .Z(n15315) );
  XOR U15158 ( .A(n15171), .B(n15317), .Z(n7638) );
  IV U15159 ( .A(n15170), .Z(n15317) );
  XNOR U15160 ( .A(n15167), .B(n15318), .Z(n15170) );
  XOR U15161 ( .A(n15319), .B(n15320), .Z(n15167) );
  ANDN U15162 ( .A(n15321), .B(n15322), .Z(n15320) );
  XNOR U15163 ( .A(n15319), .B(n15323), .Z(n15321) );
  XOR U15164 ( .A(n15178), .B(n15324), .Z(n15171) );
  IV U15165 ( .A(n15177), .Z(n15324) );
  XNOR U15166 ( .A(n15174), .B(n15325), .Z(n15177) );
  XOR U15167 ( .A(n15326), .B(n15327), .Z(n15174) );
  ANDN U15168 ( .A(n15328), .B(n15329), .Z(n15327) );
  XNOR U15169 ( .A(n15326), .B(n15330), .Z(n15328) );
  XOR U15170 ( .A(n15185), .B(n15331), .Z(n15178) );
  IV U15171 ( .A(n15184), .Z(n15331) );
  XNOR U15172 ( .A(n15181), .B(n15332), .Z(n15184) );
  XOR U15173 ( .A(n15333), .B(n15334), .Z(n15181) );
  ANDN U15174 ( .A(n15335), .B(n15336), .Z(n15334) );
  XNOR U15175 ( .A(n15333), .B(n15337), .Z(n15335) );
  XOR U15176 ( .A(n15192), .B(n15338), .Z(n15185) );
  IV U15177 ( .A(n15191), .Z(n15338) );
  XNOR U15178 ( .A(n15188), .B(n15339), .Z(n15191) );
  XOR U15179 ( .A(n15340), .B(n15341), .Z(n15188) );
  ANDN U15180 ( .A(n15342), .B(n15343), .Z(n15341) );
  XNOR U15181 ( .A(n15340), .B(n15344), .Z(n15342) );
  XOR U15182 ( .A(n15199), .B(n15345), .Z(n15192) );
  IV U15183 ( .A(n15198), .Z(n15345) );
  XNOR U15184 ( .A(n15195), .B(n15346), .Z(n15198) );
  XOR U15185 ( .A(n15347), .B(n15348), .Z(n15195) );
  ANDN U15186 ( .A(n15349), .B(n15350), .Z(n15348) );
  XNOR U15187 ( .A(n15347), .B(n15351), .Z(n15349) );
  XOR U15188 ( .A(n15206), .B(n15352), .Z(n15199) );
  IV U15189 ( .A(n15205), .Z(n15352) );
  XNOR U15190 ( .A(n15202), .B(n15353), .Z(n15205) );
  XOR U15191 ( .A(n15354), .B(n15355), .Z(n15202) );
  ANDN U15192 ( .A(n15356), .B(n15357), .Z(n15355) );
  XNOR U15193 ( .A(n15354), .B(n15358), .Z(n15356) );
  XOR U15194 ( .A(n15213), .B(n15359), .Z(n15206) );
  IV U15195 ( .A(n15212), .Z(n15359) );
  XNOR U15196 ( .A(n15209), .B(n15360), .Z(n15212) );
  XOR U15197 ( .A(n15361), .B(n15362), .Z(n15209) );
  ANDN U15198 ( .A(n15363), .B(n15364), .Z(n15362) );
  XNOR U15199 ( .A(n15361), .B(n15365), .Z(n15363) );
  XOR U15200 ( .A(n15220), .B(n15366), .Z(n15213) );
  IV U15201 ( .A(n15219), .Z(n15366) );
  XNOR U15202 ( .A(n15216), .B(n15367), .Z(n15219) );
  XOR U15203 ( .A(n15368), .B(n15369), .Z(n15216) );
  ANDN U15204 ( .A(n15370), .B(n15371), .Z(n15369) );
  XNOR U15205 ( .A(n15368), .B(n15372), .Z(n15370) );
  XOR U15206 ( .A(n15227), .B(n15373), .Z(n15220) );
  IV U15207 ( .A(n15226), .Z(n15373) );
  XNOR U15208 ( .A(n15223), .B(n15374), .Z(n15226) );
  XOR U15209 ( .A(n15375), .B(n15376), .Z(n15223) );
  ANDN U15210 ( .A(n15377), .B(n15378), .Z(n15376) );
  XNOR U15211 ( .A(n15375), .B(n15379), .Z(n15377) );
  XOR U15212 ( .A(n15234), .B(n15380), .Z(n15227) );
  IV U15213 ( .A(n15233), .Z(n15380) );
  XNOR U15214 ( .A(n15230), .B(n15381), .Z(n15233) );
  XOR U15215 ( .A(n15382), .B(n15383), .Z(n15230) );
  ANDN U15216 ( .A(n15384), .B(n15385), .Z(n15383) );
  XNOR U15217 ( .A(n15382), .B(n15386), .Z(n15384) );
  XOR U15218 ( .A(n15241), .B(n15387), .Z(n15234) );
  IV U15219 ( .A(n15240), .Z(n15387) );
  XNOR U15220 ( .A(n15237), .B(n15388), .Z(n15240) );
  XOR U15221 ( .A(n15389), .B(n15390), .Z(n15237) );
  ANDN U15222 ( .A(n15391), .B(n15392), .Z(n15390) );
  XNOR U15223 ( .A(n15389), .B(n15393), .Z(n15391) );
  XOR U15224 ( .A(n15247), .B(n15394), .Z(n15241) );
  IV U15225 ( .A(n15246), .Z(n15394) );
  XNOR U15226 ( .A(n15243), .B(n15388), .Z(n15246) );
  AND U15227 ( .A(n15553), .B(n15236), .Z(n15388) );
  XOR U15228 ( .A(n15395), .B(n15396), .Z(n15243) );
  ANDN U15229 ( .A(n15397), .B(n15398), .Z(n15396) );
  XNOR U15230 ( .A(n15395), .B(n15399), .Z(n15397) );
  XOR U15231 ( .A(n15253), .B(n15400), .Z(n15247) );
  IV U15232 ( .A(n15252), .Z(n15400) );
  XNOR U15233 ( .A(n15249), .B(n15381), .Z(n15252) );
  AND U15234 ( .A(n15896), .B(n14945), .Z(n15381) );
  XOR U15235 ( .A(n15401), .B(n15402), .Z(n15249) );
  ANDN U15236 ( .A(n15403), .B(n15404), .Z(n15402) );
  XNOR U15237 ( .A(n15401), .B(n15405), .Z(n15403) );
  XOR U15238 ( .A(n15259), .B(n15406), .Z(n15253) );
  IV U15239 ( .A(n15258), .Z(n15406) );
  XNOR U15240 ( .A(n15255), .B(n15374), .Z(n15258) );
  AND U15241 ( .A(n16265), .B(n14680), .Z(n15374) );
  XOR U15242 ( .A(n15407), .B(n15408), .Z(n15255) );
  ANDN U15243 ( .A(n15409), .B(n15410), .Z(n15408) );
  XNOR U15244 ( .A(n15407), .B(n15411), .Z(n15409) );
  XOR U15245 ( .A(n15265), .B(n15412), .Z(n15259) );
  IV U15246 ( .A(n15264), .Z(n15412) );
  XNOR U15247 ( .A(n15261), .B(n15367), .Z(n15264) );
  AND U15248 ( .A(n16657), .B(n14441), .Z(n15367) );
  XOR U15249 ( .A(n15413), .B(n15414), .Z(n15261) );
  ANDN U15250 ( .A(n15415), .B(n15416), .Z(n15414) );
  XNOR U15251 ( .A(n15413), .B(n15417), .Z(n15415) );
  XOR U15252 ( .A(n15271), .B(n15418), .Z(n15265) );
  IV U15253 ( .A(n15270), .Z(n15418) );
  XNOR U15254 ( .A(n15267), .B(n15360), .Z(n15270) );
  AND U15255 ( .A(n17567), .B(n14228), .Z(n15360) );
  XOR U15256 ( .A(n15419), .B(n15420), .Z(n15267) );
  ANDN U15257 ( .A(n15421), .B(n15422), .Z(n15420) );
  XNOR U15258 ( .A(n15419), .B(n15423), .Z(n15421) );
  XOR U15259 ( .A(n15277), .B(n15424), .Z(n15271) );
  IV U15260 ( .A(n15276), .Z(n15424) );
  XNOR U15261 ( .A(n15273), .B(n15353), .Z(n15276) );
  AND U15262 ( .A(n17688), .B(n14041), .Z(n15353) );
  XOR U15263 ( .A(n15425), .B(n15426), .Z(n15273) );
  ANDN U15264 ( .A(n15427), .B(n15428), .Z(n15426) );
  XNOR U15265 ( .A(n15425), .B(n15429), .Z(n15427) );
  XOR U15266 ( .A(n15283), .B(n15430), .Z(n15277) );
  IV U15267 ( .A(n15282), .Z(n15430) );
  XNOR U15268 ( .A(n15279), .B(n15346), .Z(n15282) );
  AND U15269 ( .A(n17814), .B(n13880), .Z(n15346) );
  XOR U15270 ( .A(n15431), .B(n15432), .Z(n15279) );
  ANDN U15271 ( .A(n15433), .B(n15434), .Z(n15432) );
  XNOR U15272 ( .A(n15431), .B(n15435), .Z(n15433) );
  XOR U15273 ( .A(n15289), .B(n15436), .Z(n15283) );
  IV U15274 ( .A(n15288), .Z(n15436) );
  XNOR U15275 ( .A(n15285), .B(n15339), .Z(n15288) );
  AND U15276 ( .A(n17945), .B(n13745), .Z(n15339) );
  XOR U15277 ( .A(n15437), .B(n15438), .Z(n15285) );
  ANDN U15278 ( .A(n15439), .B(n15440), .Z(n15438) );
  XNOR U15279 ( .A(n15437), .B(n15441), .Z(n15439) );
  XOR U15280 ( .A(n15295), .B(n15442), .Z(n15289) );
  IV U15281 ( .A(n15294), .Z(n15442) );
  XNOR U15282 ( .A(n15291), .B(n15332), .Z(n15294) );
  AND U15283 ( .A(n18081), .B(n13636), .Z(n15332) );
  XOR U15284 ( .A(n15443), .B(n15444), .Z(n15291) );
  ANDN U15285 ( .A(n15445), .B(n15446), .Z(n15444) );
  XNOR U15286 ( .A(n15443), .B(n15447), .Z(n15445) );
  XOR U15287 ( .A(n15301), .B(n15448), .Z(n15295) );
  IV U15288 ( .A(n15300), .Z(n15448) );
  XNOR U15289 ( .A(n15297), .B(n15325), .Z(n15300) );
  AND U15290 ( .A(n18222), .B(n13553), .Z(n15325) );
  XOR U15291 ( .A(n15449), .B(n15450), .Z(n15297) );
  ANDN U15292 ( .A(n15451), .B(n15452), .Z(n15450) );
  XNOR U15293 ( .A(n15449), .B(n15453), .Z(n15451) );
  XOR U15294 ( .A(n15307), .B(n15454), .Z(n15301) );
  IV U15295 ( .A(n15306), .Z(n15454) );
  XNOR U15296 ( .A(n15303), .B(n15318), .Z(n15306) );
  AND U15297 ( .A(n18368), .B(n13496), .Z(n15318) );
  XOR U15298 ( .A(n15455), .B(n15456), .Z(n15303) );
  ANDN U15299 ( .A(n15457), .B(n15458), .Z(n15456) );
  XNOR U15300 ( .A(n15455), .B(n15459), .Z(n15457) );
  XOR U15301 ( .A(n15312), .B(n15460), .Z(n15307) );
  IV U15302 ( .A(n15311), .Z(n15460) );
  XNOR U15303 ( .A(n15308), .B(n15316), .Z(n15311) );
  AND U15304 ( .A(n13470), .B(n18519), .Z(n15316) );
  XOR U15305 ( .A(n15461), .B(n15462), .Z(n15308) );
  ANDN U15306 ( .A(n15463), .B(n15464), .Z(n15462) );
  XNOR U15307 ( .A(n15461), .B(n15465), .Z(n15463) );
  XNOR U15308 ( .A(n15466), .B(n15467), .Z(n15312) );
  ANDN U15309 ( .A(n15468), .B(n15469), .Z(n15467) );
  XNOR U15310 ( .A(n15466), .B(n15470), .Z(n15468) );
  XOR U15311 ( .A(n15471), .B(n15472), .Z(n15313) );
  ANDN U15312 ( .A(n15473), .B(n7898), .Z(n15472) );
  XNOR U15313 ( .A(n15471), .B(n15474), .Z(n7898) );
  XNOR U15314 ( .A(n15471), .B(n7896), .Z(n15473) );
  XOR U15315 ( .A(n15323), .B(n15475), .Z(n7896) );
  IV U15316 ( .A(n15322), .Z(n15475) );
  XNOR U15317 ( .A(n15319), .B(n15476), .Z(n15322) );
  XOR U15318 ( .A(n15477), .B(n15478), .Z(n15319) );
  ANDN U15319 ( .A(n15479), .B(n15480), .Z(n15478) );
  XNOR U15320 ( .A(n15477), .B(n15481), .Z(n15479) );
  XOR U15321 ( .A(n15330), .B(n15482), .Z(n15323) );
  IV U15322 ( .A(n15329), .Z(n15482) );
  XNOR U15323 ( .A(n15326), .B(n15483), .Z(n15329) );
  XOR U15324 ( .A(n15484), .B(n15485), .Z(n15326) );
  ANDN U15325 ( .A(n15486), .B(n15487), .Z(n15485) );
  XNOR U15326 ( .A(n15484), .B(n15488), .Z(n15486) );
  XOR U15327 ( .A(n15337), .B(n15489), .Z(n15330) );
  IV U15328 ( .A(n15336), .Z(n15489) );
  XNOR U15329 ( .A(n15333), .B(n15490), .Z(n15336) );
  XOR U15330 ( .A(n15491), .B(n15492), .Z(n15333) );
  ANDN U15331 ( .A(n15493), .B(n15494), .Z(n15492) );
  XNOR U15332 ( .A(n15491), .B(n15495), .Z(n15493) );
  XOR U15333 ( .A(n15344), .B(n15496), .Z(n15337) );
  IV U15334 ( .A(n15343), .Z(n15496) );
  XNOR U15335 ( .A(n15340), .B(n15497), .Z(n15343) );
  XOR U15336 ( .A(n15498), .B(n15499), .Z(n15340) );
  ANDN U15337 ( .A(n15500), .B(n15501), .Z(n15499) );
  XNOR U15338 ( .A(n15498), .B(n15502), .Z(n15500) );
  XOR U15339 ( .A(n15351), .B(n15503), .Z(n15344) );
  IV U15340 ( .A(n15350), .Z(n15503) );
  XNOR U15341 ( .A(n15347), .B(n15504), .Z(n15350) );
  XOR U15342 ( .A(n15505), .B(n15506), .Z(n15347) );
  ANDN U15343 ( .A(n15507), .B(n15508), .Z(n15506) );
  XNOR U15344 ( .A(n15505), .B(n15509), .Z(n15507) );
  XOR U15345 ( .A(n15358), .B(n15510), .Z(n15351) );
  IV U15346 ( .A(n15357), .Z(n15510) );
  XNOR U15347 ( .A(n15354), .B(n15511), .Z(n15357) );
  XOR U15348 ( .A(n15512), .B(n15513), .Z(n15354) );
  ANDN U15349 ( .A(n15514), .B(n15515), .Z(n15513) );
  XNOR U15350 ( .A(n15512), .B(n15516), .Z(n15514) );
  XOR U15351 ( .A(n15365), .B(n15517), .Z(n15358) );
  IV U15352 ( .A(n15364), .Z(n15517) );
  XNOR U15353 ( .A(n15361), .B(n15518), .Z(n15364) );
  XOR U15354 ( .A(n15519), .B(n15520), .Z(n15361) );
  ANDN U15355 ( .A(n15521), .B(n15522), .Z(n15520) );
  XNOR U15356 ( .A(n15519), .B(n15523), .Z(n15521) );
  XOR U15357 ( .A(n15372), .B(n15524), .Z(n15365) );
  IV U15358 ( .A(n15371), .Z(n15524) );
  XNOR U15359 ( .A(n15368), .B(n15525), .Z(n15371) );
  XOR U15360 ( .A(n15526), .B(n15527), .Z(n15368) );
  ANDN U15361 ( .A(n15528), .B(n15529), .Z(n15527) );
  XNOR U15362 ( .A(n15526), .B(n15530), .Z(n15528) );
  XOR U15363 ( .A(n15379), .B(n15531), .Z(n15372) );
  IV U15364 ( .A(n15378), .Z(n15531) );
  XNOR U15365 ( .A(n15375), .B(n15532), .Z(n15378) );
  XOR U15366 ( .A(n15533), .B(n15534), .Z(n15375) );
  ANDN U15367 ( .A(n15535), .B(n15536), .Z(n15534) );
  XNOR U15368 ( .A(n15533), .B(n15537), .Z(n15535) );
  XOR U15369 ( .A(n15386), .B(n15538), .Z(n15379) );
  IV U15370 ( .A(n15385), .Z(n15538) );
  XNOR U15371 ( .A(n15382), .B(n15539), .Z(n15385) );
  XOR U15372 ( .A(n15540), .B(n15541), .Z(n15382) );
  ANDN U15373 ( .A(n15542), .B(n15543), .Z(n15541) );
  XNOR U15374 ( .A(n15540), .B(n15544), .Z(n15542) );
  XOR U15375 ( .A(n15393), .B(n15545), .Z(n15386) );
  IV U15376 ( .A(n15392), .Z(n15545) );
  XNOR U15377 ( .A(n15389), .B(n15546), .Z(n15392) );
  XOR U15378 ( .A(n15547), .B(n15548), .Z(n15389) );
  ANDN U15379 ( .A(n15549), .B(n15550), .Z(n15548) );
  XNOR U15380 ( .A(n15547), .B(n15551), .Z(n15549) );
  XOR U15381 ( .A(n15399), .B(n15552), .Z(n15393) );
  IV U15382 ( .A(n15398), .Z(n15552) );
  XNOR U15383 ( .A(n15395), .B(n15553), .Z(n15398) );
  XOR U15384 ( .A(n15554), .B(n15555), .Z(n15395) );
  ANDN U15385 ( .A(n15556), .B(n15557), .Z(n15555) );
  XNOR U15386 ( .A(n15554), .B(n15558), .Z(n15556) );
  XOR U15387 ( .A(n15405), .B(n15559), .Z(n15399) );
  IV U15388 ( .A(n15404), .Z(n15559) );
  XNOR U15389 ( .A(n15401), .B(n15546), .Z(n15404) );
  AND U15390 ( .A(n15896), .B(n15236), .Z(n15546) );
  XOR U15391 ( .A(n15560), .B(n15561), .Z(n15401) );
  ANDN U15392 ( .A(n15562), .B(n15563), .Z(n15561) );
  XNOR U15393 ( .A(n15560), .B(n15564), .Z(n15562) );
  XOR U15394 ( .A(n15411), .B(n15565), .Z(n15405) );
  IV U15395 ( .A(n15410), .Z(n15565) );
  XNOR U15396 ( .A(n15407), .B(n15539), .Z(n15410) );
  AND U15397 ( .A(n16265), .B(n14945), .Z(n15539) );
  XOR U15398 ( .A(n15566), .B(n15567), .Z(n15407) );
  ANDN U15399 ( .A(n15568), .B(n15569), .Z(n15567) );
  XNOR U15400 ( .A(n15566), .B(n15570), .Z(n15568) );
  XOR U15401 ( .A(n15417), .B(n15571), .Z(n15411) );
  IV U15402 ( .A(n15416), .Z(n15571) );
  XNOR U15403 ( .A(n15413), .B(n15532), .Z(n15416) );
  AND U15404 ( .A(n16657), .B(n14680), .Z(n15532) );
  XOR U15405 ( .A(n15572), .B(n15573), .Z(n15413) );
  ANDN U15406 ( .A(n15574), .B(n15575), .Z(n15573) );
  XNOR U15407 ( .A(n15572), .B(n15576), .Z(n15574) );
  XOR U15408 ( .A(n15423), .B(n15577), .Z(n15417) );
  IV U15409 ( .A(n15422), .Z(n15577) );
  XNOR U15410 ( .A(n15419), .B(n15525), .Z(n15422) );
  AND U15411 ( .A(n17567), .B(n14441), .Z(n15525) );
  XOR U15412 ( .A(n15578), .B(n15579), .Z(n15419) );
  ANDN U15413 ( .A(n15580), .B(n15581), .Z(n15579) );
  XNOR U15414 ( .A(n15578), .B(n15582), .Z(n15580) );
  XOR U15415 ( .A(n15429), .B(n15583), .Z(n15423) );
  IV U15416 ( .A(n15428), .Z(n15583) );
  XNOR U15417 ( .A(n15425), .B(n15518), .Z(n15428) );
  AND U15418 ( .A(n17688), .B(n14228), .Z(n15518) );
  XOR U15419 ( .A(n15584), .B(n15585), .Z(n15425) );
  ANDN U15420 ( .A(n15586), .B(n15587), .Z(n15585) );
  XNOR U15421 ( .A(n15584), .B(n15588), .Z(n15586) );
  XOR U15422 ( .A(n15435), .B(n15589), .Z(n15429) );
  IV U15423 ( .A(n15434), .Z(n15589) );
  XNOR U15424 ( .A(n15431), .B(n15511), .Z(n15434) );
  AND U15425 ( .A(n17814), .B(n14041), .Z(n15511) );
  XOR U15426 ( .A(n15590), .B(n15591), .Z(n15431) );
  ANDN U15427 ( .A(n15592), .B(n15593), .Z(n15591) );
  XNOR U15428 ( .A(n15590), .B(n15594), .Z(n15592) );
  XOR U15429 ( .A(n15441), .B(n15595), .Z(n15435) );
  IV U15430 ( .A(n15440), .Z(n15595) );
  XNOR U15431 ( .A(n15437), .B(n15504), .Z(n15440) );
  AND U15432 ( .A(n17945), .B(n13880), .Z(n15504) );
  XOR U15433 ( .A(n15596), .B(n15597), .Z(n15437) );
  ANDN U15434 ( .A(n15598), .B(n15599), .Z(n15597) );
  XNOR U15435 ( .A(n15596), .B(n15600), .Z(n15598) );
  XOR U15436 ( .A(n15447), .B(n15601), .Z(n15441) );
  IV U15437 ( .A(n15446), .Z(n15601) );
  XNOR U15438 ( .A(n15443), .B(n15497), .Z(n15446) );
  AND U15439 ( .A(n18081), .B(n13745), .Z(n15497) );
  XOR U15440 ( .A(n15602), .B(n15603), .Z(n15443) );
  ANDN U15441 ( .A(n15604), .B(n15605), .Z(n15603) );
  XNOR U15442 ( .A(n15602), .B(n15606), .Z(n15604) );
  XOR U15443 ( .A(n15453), .B(n15607), .Z(n15447) );
  IV U15444 ( .A(n15452), .Z(n15607) );
  XNOR U15445 ( .A(n15449), .B(n15490), .Z(n15452) );
  AND U15446 ( .A(n18222), .B(n13636), .Z(n15490) );
  XOR U15447 ( .A(n15608), .B(n15609), .Z(n15449) );
  ANDN U15448 ( .A(n15610), .B(n15611), .Z(n15609) );
  XNOR U15449 ( .A(n15608), .B(n15612), .Z(n15610) );
  XOR U15450 ( .A(n15459), .B(n15613), .Z(n15453) );
  IV U15451 ( .A(n15458), .Z(n15613) );
  XNOR U15452 ( .A(n15455), .B(n15483), .Z(n15458) );
  AND U15453 ( .A(n18368), .B(n13553), .Z(n15483) );
  XOR U15454 ( .A(n15614), .B(n15615), .Z(n15455) );
  ANDN U15455 ( .A(n15616), .B(n15617), .Z(n15615) );
  XNOR U15456 ( .A(n15614), .B(n15618), .Z(n15616) );
  XOR U15457 ( .A(n15465), .B(n15619), .Z(n15459) );
  IV U15458 ( .A(n15464), .Z(n15619) );
  XNOR U15459 ( .A(n15461), .B(n15476), .Z(n15464) );
  AND U15460 ( .A(n18519), .B(n13496), .Z(n15476) );
  XOR U15461 ( .A(n15620), .B(n15621), .Z(n15461) );
  ANDN U15462 ( .A(n15622), .B(n15623), .Z(n15621) );
  XNOR U15463 ( .A(n15620), .B(n15624), .Z(n15622) );
  XOR U15464 ( .A(n15470), .B(n15625), .Z(n15465) );
  IV U15465 ( .A(n15469), .Z(n15625) );
  XNOR U15466 ( .A(n15466), .B(n15474), .Z(n15469) );
  AND U15467 ( .A(n13470), .B(n18675), .Z(n15474) );
  XOR U15468 ( .A(n15626), .B(n15627), .Z(n15466) );
  ANDN U15469 ( .A(n15628), .B(n15629), .Z(n15627) );
  XNOR U15470 ( .A(n15626), .B(n15630), .Z(n15628) );
  XNOR U15471 ( .A(n15631), .B(n15632), .Z(n15470) );
  ANDN U15472 ( .A(n15633), .B(n15634), .Z(n15632) );
  XNOR U15473 ( .A(n15631), .B(n15635), .Z(n15633) );
  XOR U15474 ( .A(n15636), .B(n15637), .Z(n15471) );
  ANDN U15475 ( .A(n15638), .B(n8149), .Z(n15637) );
  XNOR U15476 ( .A(n15636), .B(n15639), .Z(n8149) );
  XNOR U15477 ( .A(n15636), .B(n8147), .Z(n15638) );
  XOR U15478 ( .A(n15481), .B(n15640), .Z(n8147) );
  IV U15479 ( .A(n15480), .Z(n15640) );
  XNOR U15480 ( .A(n15477), .B(n15641), .Z(n15480) );
  XOR U15481 ( .A(n15642), .B(n15643), .Z(n15477) );
  ANDN U15482 ( .A(n15644), .B(n15645), .Z(n15643) );
  XNOR U15483 ( .A(n15642), .B(n15646), .Z(n15644) );
  XOR U15484 ( .A(n15488), .B(n15647), .Z(n15481) );
  IV U15485 ( .A(n15487), .Z(n15647) );
  XNOR U15486 ( .A(n15484), .B(n15648), .Z(n15487) );
  XOR U15487 ( .A(n15649), .B(n15650), .Z(n15484) );
  ANDN U15488 ( .A(n15651), .B(n15652), .Z(n15650) );
  XNOR U15489 ( .A(n15649), .B(n15653), .Z(n15651) );
  XOR U15490 ( .A(n15495), .B(n15654), .Z(n15488) );
  IV U15491 ( .A(n15494), .Z(n15654) );
  XNOR U15492 ( .A(n15491), .B(n15655), .Z(n15494) );
  XOR U15493 ( .A(n15656), .B(n15657), .Z(n15491) );
  ANDN U15494 ( .A(n15658), .B(n15659), .Z(n15657) );
  XNOR U15495 ( .A(n15656), .B(n15660), .Z(n15658) );
  XOR U15496 ( .A(n15502), .B(n15661), .Z(n15495) );
  IV U15497 ( .A(n15501), .Z(n15661) );
  XNOR U15498 ( .A(n15498), .B(n15662), .Z(n15501) );
  XOR U15499 ( .A(n15663), .B(n15664), .Z(n15498) );
  ANDN U15500 ( .A(n15665), .B(n15666), .Z(n15664) );
  XNOR U15501 ( .A(n15663), .B(n15667), .Z(n15665) );
  XOR U15502 ( .A(n15509), .B(n15668), .Z(n15502) );
  IV U15503 ( .A(n15508), .Z(n15668) );
  XNOR U15504 ( .A(n15505), .B(n15669), .Z(n15508) );
  XOR U15505 ( .A(n15670), .B(n15671), .Z(n15505) );
  ANDN U15506 ( .A(n15672), .B(n15673), .Z(n15671) );
  XNOR U15507 ( .A(n15670), .B(n15674), .Z(n15672) );
  XOR U15508 ( .A(n15516), .B(n15675), .Z(n15509) );
  IV U15509 ( .A(n15515), .Z(n15675) );
  XNOR U15510 ( .A(n15512), .B(n15676), .Z(n15515) );
  XOR U15511 ( .A(n15677), .B(n15678), .Z(n15512) );
  ANDN U15512 ( .A(n15679), .B(n15680), .Z(n15678) );
  XNOR U15513 ( .A(n15677), .B(n15681), .Z(n15679) );
  XOR U15514 ( .A(n15523), .B(n15682), .Z(n15516) );
  IV U15515 ( .A(n15522), .Z(n15682) );
  XNOR U15516 ( .A(n15519), .B(n15683), .Z(n15522) );
  XOR U15517 ( .A(n15684), .B(n15685), .Z(n15519) );
  ANDN U15518 ( .A(n15686), .B(n15687), .Z(n15685) );
  XNOR U15519 ( .A(n15684), .B(n15688), .Z(n15686) );
  XOR U15520 ( .A(n15530), .B(n15689), .Z(n15523) );
  IV U15521 ( .A(n15529), .Z(n15689) );
  XNOR U15522 ( .A(n15526), .B(n15690), .Z(n15529) );
  XOR U15523 ( .A(n15691), .B(n15692), .Z(n15526) );
  ANDN U15524 ( .A(n15693), .B(n15694), .Z(n15692) );
  XNOR U15525 ( .A(n15691), .B(n15695), .Z(n15693) );
  XOR U15526 ( .A(n15537), .B(n15696), .Z(n15530) );
  IV U15527 ( .A(n15536), .Z(n15696) );
  XNOR U15528 ( .A(n15533), .B(n15697), .Z(n15536) );
  XOR U15529 ( .A(n15698), .B(n15699), .Z(n15533) );
  ANDN U15530 ( .A(n15700), .B(n15701), .Z(n15699) );
  XNOR U15531 ( .A(n15698), .B(n15702), .Z(n15700) );
  XOR U15532 ( .A(n15544), .B(n15703), .Z(n15537) );
  IV U15533 ( .A(n15543), .Z(n15703) );
  XNOR U15534 ( .A(n15540), .B(n15704), .Z(n15543) );
  XOR U15535 ( .A(n15705), .B(n15706), .Z(n15540) );
  ANDN U15536 ( .A(n15707), .B(n15708), .Z(n15706) );
  XNOR U15537 ( .A(n15705), .B(n15709), .Z(n15707) );
  XOR U15538 ( .A(n15551), .B(n15710), .Z(n15544) );
  IV U15539 ( .A(n15550), .Z(n15710) );
  XNOR U15540 ( .A(n15547), .B(n15711), .Z(n15550) );
  XOR U15541 ( .A(n15712), .B(n15713), .Z(n15547) );
  ANDN U15542 ( .A(n15714), .B(n15715), .Z(n15713) );
  XNOR U15543 ( .A(n15712), .B(n15716), .Z(n15714) );
  XOR U15544 ( .A(n15558), .B(n15717), .Z(n15551) );
  IV U15545 ( .A(n15557), .Z(n15717) );
  XNOR U15546 ( .A(n15554), .B(n15718), .Z(n15557) );
  XOR U15547 ( .A(n15719), .B(n15720), .Z(n15554) );
  ANDN U15548 ( .A(n15721), .B(n15722), .Z(n15720) );
  XNOR U15549 ( .A(n15719), .B(n15723), .Z(n15721) );
  XOR U15550 ( .A(n15564), .B(n15724), .Z(n15558) );
  IV U15551 ( .A(n15563), .Z(n15724) );
  XNOR U15552 ( .A(n15560), .B(n15718), .Z(n15563) );
  AND U15553 ( .A(n15896), .B(n15553), .Z(n15718) );
  XOR U15554 ( .A(n15725), .B(n15726), .Z(n15560) );
  ANDN U15555 ( .A(n15727), .B(n15728), .Z(n15726) );
  XNOR U15556 ( .A(n15725), .B(n15729), .Z(n15727) );
  XOR U15557 ( .A(n15570), .B(n15730), .Z(n15564) );
  IV U15558 ( .A(n15569), .Z(n15730) );
  XNOR U15559 ( .A(n15566), .B(n15711), .Z(n15569) );
  AND U15560 ( .A(n16265), .B(n15236), .Z(n15711) );
  XOR U15561 ( .A(n15731), .B(n15732), .Z(n15566) );
  ANDN U15562 ( .A(n15733), .B(n15734), .Z(n15732) );
  XNOR U15563 ( .A(n15731), .B(n15735), .Z(n15733) );
  XOR U15564 ( .A(n15576), .B(n15736), .Z(n15570) );
  IV U15565 ( .A(n15575), .Z(n15736) );
  XNOR U15566 ( .A(n15572), .B(n15704), .Z(n15575) );
  AND U15567 ( .A(n16657), .B(n14945), .Z(n15704) );
  XOR U15568 ( .A(n15737), .B(n15738), .Z(n15572) );
  ANDN U15569 ( .A(n15739), .B(n15740), .Z(n15738) );
  XNOR U15570 ( .A(n15737), .B(n15741), .Z(n15739) );
  XOR U15571 ( .A(n15582), .B(n15742), .Z(n15576) );
  IV U15572 ( .A(n15581), .Z(n15742) );
  XNOR U15573 ( .A(n15578), .B(n15697), .Z(n15581) );
  AND U15574 ( .A(n17567), .B(n14680), .Z(n15697) );
  XOR U15575 ( .A(n15743), .B(n15744), .Z(n15578) );
  ANDN U15576 ( .A(n15745), .B(n15746), .Z(n15744) );
  XNOR U15577 ( .A(n15743), .B(n15747), .Z(n15745) );
  XOR U15578 ( .A(n15588), .B(n15748), .Z(n15582) );
  IV U15579 ( .A(n15587), .Z(n15748) );
  XNOR U15580 ( .A(n15584), .B(n15690), .Z(n15587) );
  AND U15581 ( .A(n17688), .B(n14441), .Z(n15690) );
  XOR U15582 ( .A(n15749), .B(n15750), .Z(n15584) );
  ANDN U15583 ( .A(n15751), .B(n15752), .Z(n15750) );
  XNOR U15584 ( .A(n15749), .B(n15753), .Z(n15751) );
  XOR U15585 ( .A(n15594), .B(n15754), .Z(n15588) );
  IV U15586 ( .A(n15593), .Z(n15754) );
  XNOR U15587 ( .A(n15590), .B(n15683), .Z(n15593) );
  AND U15588 ( .A(n17814), .B(n14228), .Z(n15683) );
  XOR U15589 ( .A(n15755), .B(n15756), .Z(n15590) );
  ANDN U15590 ( .A(n15757), .B(n15758), .Z(n15756) );
  XNOR U15591 ( .A(n15755), .B(n15759), .Z(n15757) );
  XOR U15592 ( .A(n15600), .B(n15760), .Z(n15594) );
  IV U15593 ( .A(n15599), .Z(n15760) );
  XNOR U15594 ( .A(n15596), .B(n15676), .Z(n15599) );
  AND U15595 ( .A(n17945), .B(n14041), .Z(n15676) );
  XOR U15596 ( .A(n15761), .B(n15762), .Z(n15596) );
  ANDN U15597 ( .A(n15763), .B(n15764), .Z(n15762) );
  XNOR U15598 ( .A(n15761), .B(n15765), .Z(n15763) );
  XOR U15599 ( .A(n15606), .B(n15766), .Z(n15600) );
  IV U15600 ( .A(n15605), .Z(n15766) );
  XNOR U15601 ( .A(n15602), .B(n15669), .Z(n15605) );
  AND U15602 ( .A(n18081), .B(n13880), .Z(n15669) );
  XOR U15603 ( .A(n15767), .B(n15768), .Z(n15602) );
  ANDN U15604 ( .A(n15769), .B(n15770), .Z(n15768) );
  XNOR U15605 ( .A(n15767), .B(n15771), .Z(n15769) );
  XOR U15606 ( .A(n15612), .B(n15772), .Z(n15606) );
  IV U15607 ( .A(n15611), .Z(n15772) );
  XNOR U15608 ( .A(n15608), .B(n15662), .Z(n15611) );
  AND U15609 ( .A(n18222), .B(n13745), .Z(n15662) );
  XOR U15610 ( .A(n15773), .B(n15774), .Z(n15608) );
  ANDN U15611 ( .A(n15775), .B(n15776), .Z(n15774) );
  XNOR U15612 ( .A(n15773), .B(n15777), .Z(n15775) );
  XOR U15613 ( .A(n15618), .B(n15778), .Z(n15612) );
  IV U15614 ( .A(n15617), .Z(n15778) );
  XNOR U15615 ( .A(n15614), .B(n15655), .Z(n15617) );
  AND U15616 ( .A(n18368), .B(n13636), .Z(n15655) );
  XOR U15617 ( .A(n15779), .B(n15780), .Z(n15614) );
  ANDN U15618 ( .A(n15781), .B(n15782), .Z(n15780) );
  XNOR U15619 ( .A(n15779), .B(n15783), .Z(n15781) );
  XOR U15620 ( .A(n15624), .B(n15784), .Z(n15618) );
  IV U15621 ( .A(n15623), .Z(n15784) );
  XNOR U15622 ( .A(n15620), .B(n15648), .Z(n15623) );
  AND U15623 ( .A(n18519), .B(n13553), .Z(n15648) );
  XOR U15624 ( .A(n15785), .B(n15786), .Z(n15620) );
  ANDN U15625 ( .A(n15787), .B(n15788), .Z(n15786) );
  XNOR U15626 ( .A(n15785), .B(n15789), .Z(n15787) );
  XOR U15627 ( .A(n15630), .B(n15790), .Z(n15624) );
  IV U15628 ( .A(n15629), .Z(n15790) );
  XNOR U15629 ( .A(n15626), .B(n15641), .Z(n15629) );
  AND U15630 ( .A(n18675), .B(n13496), .Z(n15641) );
  XOR U15631 ( .A(n15791), .B(n15792), .Z(n15626) );
  ANDN U15632 ( .A(n15793), .B(n15794), .Z(n15792) );
  XNOR U15633 ( .A(n15791), .B(n15795), .Z(n15793) );
  XOR U15634 ( .A(n15635), .B(n15796), .Z(n15630) );
  IV U15635 ( .A(n15634), .Z(n15796) );
  XNOR U15636 ( .A(n15631), .B(n15639), .Z(n15634) );
  AND U15637 ( .A(n13470), .B(n18836), .Z(n15639) );
  XOR U15638 ( .A(n15797), .B(n15798), .Z(n15631) );
  ANDN U15639 ( .A(n15799), .B(n15800), .Z(n15798) );
  XNOR U15640 ( .A(n15797), .B(n15801), .Z(n15799) );
  XNOR U15641 ( .A(n15802), .B(n15803), .Z(n15635) );
  ANDN U15642 ( .A(n15804), .B(n15805), .Z(n15803) );
  XNOR U15643 ( .A(n15802), .B(n15806), .Z(n15804) );
  XOR U15644 ( .A(n15807), .B(n15808), .Z(n15636) );
  ANDN U15645 ( .A(n15809), .B(n8394), .Z(n15808) );
  XNOR U15646 ( .A(n15807), .B(n15810), .Z(n8394) );
  XNOR U15647 ( .A(n15807), .B(n8392), .Z(n15809) );
  XOR U15648 ( .A(n15646), .B(n15811), .Z(n8392) );
  IV U15649 ( .A(n15645), .Z(n15811) );
  XNOR U15650 ( .A(n15642), .B(n15812), .Z(n15645) );
  XOR U15651 ( .A(n15813), .B(n15814), .Z(n15642) );
  ANDN U15652 ( .A(n15815), .B(n15816), .Z(n15814) );
  XNOR U15653 ( .A(n15813), .B(n15817), .Z(n15815) );
  XOR U15654 ( .A(n15653), .B(n15818), .Z(n15646) );
  IV U15655 ( .A(n15652), .Z(n15818) );
  XNOR U15656 ( .A(n15649), .B(n15819), .Z(n15652) );
  XOR U15657 ( .A(n15820), .B(n15821), .Z(n15649) );
  ANDN U15658 ( .A(n15822), .B(n15823), .Z(n15821) );
  XNOR U15659 ( .A(n15820), .B(n15824), .Z(n15822) );
  XOR U15660 ( .A(n15660), .B(n15825), .Z(n15653) );
  IV U15661 ( .A(n15659), .Z(n15825) );
  XNOR U15662 ( .A(n15656), .B(n15826), .Z(n15659) );
  XOR U15663 ( .A(n15827), .B(n15828), .Z(n15656) );
  ANDN U15664 ( .A(n15829), .B(n15830), .Z(n15828) );
  XNOR U15665 ( .A(n15827), .B(n15831), .Z(n15829) );
  XOR U15666 ( .A(n15667), .B(n15832), .Z(n15660) );
  IV U15667 ( .A(n15666), .Z(n15832) );
  XNOR U15668 ( .A(n15663), .B(n15833), .Z(n15666) );
  XOR U15669 ( .A(n15834), .B(n15835), .Z(n15663) );
  ANDN U15670 ( .A(n15836), .B(n15837), .Z(n15835) );
  XNOR U15671 ( .A(n15834), .B(n15838), .Z(n15836) );
  XOR U15672 ( .A(n15674), .B(n15839), .Z(n15667) );
  IV U15673 ( .A(n15673), .Z(n15839) );
  XNOR U15674 ( .A(n15670), .B(n15840), .Z(n15673) );
  XOR U15675 ( .A(n15841), .B(n15842), .Z(n15670) );
  ANDN U15676 ( .A(n15843), .B(n15844), .Z(n15842) );
  XNOR U15677 ( .A(n15841), .B(n15845), .Z(n15843) );
  XOR U15678 ( .A(n15681), .B(n15846), .Z(n15674) );
  IV U15679 ( .A(n15680), .Z(n15846) );
  XNOR U15680 ( .A(n15677), .B(n15847), .Z(n15680) );
  XOR U15681 ( .A(n15848), .B(n15849), .Z(n15677) );
  ANDN U15682 ( .A(n15850), .B(n15851), .Z(n15849) );
  XNOR U15683 ( .A(n15848), .B(n15852), .Z(n15850) );
  XOR U15684 ( .A(n15688), .B(n15853), .Z(n15681) );
  IV U15685 ( .A(n15687), .Z(n15853) );
  XNOR U15686 ( .A(n15684), .B(n15854), .Z(n15687) );
  XOR U15687 ( .A(n15855), .B(n15856), .Z(n15684) );
  ANDN U15688 ( .A(n15857), .B(n15858), .Z(n15856) );
  XNOR U15689 ( .A(n15855), .B(n15859), .Z(n15857) );
  XOR U15690 ( .A(n15695), .B(n15860), .Z(n15688) );
  IV U15691 ( .A(n15694), .Z(n15860) );
  XNOR U15692 ( .A(n15691), .B(n15861), .Z(n15694) );
  XOR U15693 ( .A(n15862), .B(n15863), .Z(n15691) );
  ANDN U15694 ( .A(n15864), .B(n15865), .Z(n15863) );
  XNOR U15695 ( .A(n15862), .B(n15866), .Z(n15864) );
  XOR U15696 ( .A(n15702), .B(n15867), .Z(n15695) );
  IV U15697 ( .A(n15701), .Z(n15867) );
  XNOR U15698 ( .A(n15698), .B(n15868), .Z(n15701) );
  XOR U15699 ( .A(n15869), .B(n15870), .Z(n15698) );
  ANDN U15700 ( .A(n15871), .B(n15872), .Z(n15870) );
  XNOR U15701 ( .A(n15869), .B(n15873), .Z(n15871) );
  XOR U15702 ( .A(n15709), .B(n15874), .Z(n15702) );
  IV U15703 ( .A(n15708), .Z(n15874) );
  XNOR U15704 ( .A(n15705), .B(n15875), .Z(n15708) );
  XOR U15705 ( .A(n15876), .B(n15877), .Z(n15705) );
  ANDN U15706 ( .A(n15878), .B(n15879), .Z(n15877) );
  XNOR U15707 ( .A(n15876), .B(n15880), .Z(n15878) );
  XOR U15708 ( .A(n15716), .B(n15881), .Z(n15709) );
  IV U15709 ( .A(n15715), .Z(n15881) );
  XNOR U15710 ( .A(n15712), .B(n15882), .Z(n15715) );
  XOR U15711 ( .A(n15883), .B(n15884), .Z(n15712) );
  ANDN U15712 ( .A(n15885), .B(n15886), .Z(n15884) );
  XNOR U15713 ( .A(n15883), .B(n15887), .Z(n15885) );
  XOR U15714 ( .A(n15723), .B(n15888), .Z(n15716) );
  IV U15715 ( .A(n15722), .Z(n15888) );
  XNOR U15716 ( .A(n15719), .B(n15889), .Z(n15722) );
  XOR U15717 ( .A(n15890), .B(n15891), .Z(n15719) );
  ANDN U15718 ( .A(n15892), .B(n15893), .Z(n15891) );
  XNOR U15719 ( .A(n15890), .B(n15894), .Z(n15892) );
  XOR U15720 ( .A(n15729), .B(n15895), .Z(n15723) );
  IV U15721 ( .A(n15728), .Z(n15895) );
  XNOR U15722 ( .A(n15725), .B(n15896), .Z(n15728) );
  XOR U15723 ( .A(n15897), .B(n15898), .Z(n15725) );
  ANDN U15724 ( .A(n15899), .B(n15900), .Z(n15898) );
  XNOR U15725 ( .A(n15897), .B(n15901), .Z(n15899) );
  XOR U15726 ( .A(n15735), .B(n15902), .Z(n15729) );
  IV U15727 ( .A(n15734), .Z(n15902) );
  XNOR U15728 ( .A(n15731), .B(n15889), .Z(n15734) );
  AND U15729 ( .A(n16265), .B(n15553), .Z(n15889) );
  XOR U15730 ( .A(n15903), .B(n15904), .Z(n15731) );
  ANDN U15731 ( .A(n15905), .B(n15906), .Z(n15904) );
  XNOR U15732 ( .A(n15903), .B(n15907), .Z(n15905) );
  XOR U15733 ( .A(n15741), .B(n15908), .Z(n15735) );
  IV U15734 ( .A(n15740), .Z(n15908) );
  XNOR U15735 ( .A(n15737), .B(n15882), .Z(n15740) );
  AND U15736 ( .A(n16657), .B(n15236), .Z(n15882) );
  XOR U15737 ( .A(n15909), .B(n15910), .Z(n15737) );
  ANDN U15738 ( .A(n15911), .B(n15912), .Z(n15910) );
  XNOR U15739 ( .A(n15909), .B(n15913), .Z(n15911) );
  XOR U15740 ( .A(n15747), .B(n15914), .Z(n15741) );
  IV U15741 ( .A(n15746), .Z(n15914) );
  XNOR U15742 ( .A(n15743), .B(n15875), .Z(n15746) );
  AND U15743 ( .A(n17567), .B(n14945), .Z(n15875) );
  XOR U15744 ( .A(n15915), .B(n15916), .Z(n15743) );
  ANDN U15745 ( .A(n15917), .B(n15918), .Z(n15916) );
  XNOR U15746 ( .A(n15915), .B(n15919), .Z(n15917) );
  XOR U15747 ( .A(n15753), .B(n15920), .Z(n15747) );
  IV U15748 ( .A(n15752), .Z(n15920) );
  XNOR U15749 ( .A(n15749), .B(n15868), .Z(n15752) );
  AND U15750 ( .A(n17688), .B(n14680), .Z(n15868) );
  XOR U15751 ( .A(n15921), .B(n15922), .Z(n15749) );
  ANDN U15752 ( .A(n15923), .B(n15924), .Z(n15922) );
  XNOR U15753 ( .A(n15921), .B(n15925), .Z(n15923) );
  XOR U15754 ( .A(n15759), .B(n15926), .Z(n15753) );
  IV U15755 ( .A(n15758), .Z(n15926) );
  XNOR U15756 ( .A(n15755), .B(n15861), .Z(n15758) );
  AND U15757 ( .A(n17814), .B(n14441), .Z(n15861) );
  XOR U15758 ( .A(n15927), .B(n15928), .Z(n15755) );
  ANDN U15759 ( .A(n15929), .B(n15930), .Z(n15928) );
  XNOR U15760 ( .A(n15927), .B(n15931), .Z(n15929) );
  XOR U15761 ( .A(n15765), .B(n15932), .Z(n15759) );
  IV U15762 ( .A(n15764), .Z(n15932) );
  XNOR U15763 ( .A(n15761), .B(n15854), .Z(n15764) );
  AND U15764 ( .A(n17945), .B(n14228), .Z(n15854) );
  XOR U15765 ( .A(n15933), .B(n15934), .Z(n15761) );
  ANDN U15766 ( .A(n15935), .B(n15936), .Z(n15934) );
  XNOR U15767 ( .A(n15933), .B(n15937), .Z(n15935) );
  XOR U15768 ( .A(n15771), .B(n15938), .Z(n15765) );
  IV U15769 ( .A(n15770), .Z(n15938) );
  XNOR U15770 ( .A(n15767), .B(n15847), .Z(n15770) );
  AND U15771 ( .A(n18081), .B(n14041), .Z(n15847) );
  XOR U15772 ( .A(n15939), .B(n15940), .Z(n15767) );
  ANDN U15773 ( .A(n15941), .B(n15942), .Z(n15940) );
  XNOR U15774 ( .A(n15939), .B(n15943), .Z(n15941) );
  XOR U15775 ( .A(n15777), .B(n15944), .Z(n15771) );
  IV U15776 ( .A(n15776), .Z(n15944) );
  XNOR U15777 ( .A(n15773), .B(n15840), .Z(n15776) );
  AND U15778 ( .A(n18222), .B(n13880), .Z(n15840) );
  XOR U15779 ( .A(n15945), .B(n15946), .Z(n15773) );
  ANDN U15780 ( .A(n15947), .B(n15948), .Z(n15946) );
  XNOR U15781 ( .A(n15945), .B(n15949), .Z(n15947) );
  XOR U15782 ( .A(n15783), .B(n15950), .Z(n15777) );
  IV U15783 ( .A(n15782), .Z(n15950) );
  XNOR U15784 ( .A(n15779), .B(n15833), .Z(n15782) );
  AND U15785 ( .A(n18368), .B(n13745), .Z(n15833) );
  XOR U15786 ( .A(n15951), .B(n15952), .Z(n15779) );
  ANDN U15787 ( .A(n15953), .B(n15954), .Z(n15952) );
  XNOR U15788 ( .A(n15951), .B(n15955), .Z(n15953) );
  XOR U15789 ( .A(n15789), .B(n15956), .Z(n15783) );
  IV U15790 ( .A(n15788), .Z(n15956) );
  XNOR U15791 ( .A(n15785), .B(n15826), .Z(n15788) );
  AND U15792 ( .A(n18519), .B(n13636), .Z(n15826) );
  XOR U15793 ( .A(n15957), .B(n15958), .Z(n15785) );
  ANDN U15794 ( .A(n15959), .B(n15960), .Z(n15958) );
  XNOR U15795 ( .A(n15957), .B(n15961), .Z(n15959) );
  XOR U15796 ( .A(n15795), .B(n15962), .Z(n15789) );
  IV U15797 ( .A(n15794), .Z(n15962) );
  XNOR U15798 ( .A(n15791), .B(n15819), .Z(n15794) );
  AND U15799 ( .A(n18675), .B(n13553), .Z(n15819) );
  XOR U15800 ( .A(n15963), .B(n15964), .Z(n15791) );
  ANDN U15801 ( .A(n15965), .B(n15966), .Z(n15964) );
  XNOR U15802 ( .A(n15963), .B(n15967), .Z(n15965) );
  XOR U15803 ( .A(n15801), .B(n15968), .Z(n15795) );
  IV U15804 ( .A(n15800), .Z(n15968) );
  XNOR U15805 ( .A(n15797), .B(n15812), .Z(n15800) );
  AND U15806 ( .A(n18836), .B(n13496), .Z(n15812) );
  XOR U15807 ( .A(n15969), .B(n15970), .Z(n15797) );
  ANDN U15808 ( .A(n15971), .B(n15972), .Z(n15970) );
  XNOR U15809 ( .A(n15969), .B(n15973), .Z(n15971) );
  XOR U15810 ( .A(n15806), .B(n15974), .Z(n15801) );
  IV U15811 ( .A(n15805), .Z(n15974) );
  XNOR U15812 ( .A(n15802), .B(n15810), .Z(n15805) );
  AND U15813 ( .A(n13470), .B(n19002), .Z(n15810) );
  XOR U15814 ( .A(n15975), .B(n15976), .Z(n15802) );
  ANDN U15815 ( .A(n15977), .B(n15978), .Z(n15976) );
  XNOR U15816 ( .A(n15975), .B(n15979), .Z(n15977) );
  XNOR U15817 ( .A(n15980), .B(n15981), .Z(n15806) );
  ANDN U15818 ( .A(n15982), .B(n15983), .Z(n15981) );
  XNOR U15819 ( .A(n15980), .B(n15984), .Z(n15982) );
  XOR U15820 ( .A(n15985), .B(n15986), .Z(n15807) );
  ANDN U15821 ( .A(n15987), .B(n8632), .Z(n15986) );
  XNOR U15822 ( .A(n15985), .B(n15988), .Z(n8632) );
  XNOR U15823 ( .A(n15985), .B(n8630), .Z(n15987) );
  XOR U15824 ( .A(n15817), .B(n15989), .Z(n8630) );
  IV U15825 ( .A(n15816), .Z(n15989) );
  XNOR U15826 ( .A(n15813), .B(n15990), .Z(n15816) );
  XOR U15827 ( .A(n15991), .B(n15992), .Z(n15813) );
  ANDN U15828 ( .A(n15993), .B(n15994), .Z(n15992) );
  XNOR U15829 ( .A(n15991), .B(n15995), .Z(n15993) );
  XOR U15830 ( .A(n15824), .B(n15996), .Z(n15817) );
  IV U15831 ( .A(n15823), .Z(n15996) );
  XNOR U15832 ( .A(n15820), .B(n15997), .Z(n15823) );
  XOR U15833 ( .A(n15998), .B(n15999), .Z(n15820) );
  ANDN U15834 ( .A(n16000), .B(n16001), .Z(n15999) );
  XNOR U15835 ( .A(n15998), .B(n16002), .Z(n16000) );
  XOR U15836 ( .A(n15831), .B(n16003), .Z(n15824) );
  IV U15837 ( .A(n15830), .Z(n16003) );
  XNOR U15838 ( .A(n15827), .B(n16004), .Z(n15830) );
  XOR U15839 ( .A(n16005), .B(n16006), .Z(n15827) );
  ANDN U15840 ( .A(n16007), .B(n16008), .Z(n16006) );
  XNOR U15841 ( .A(n16005), .B(n16009), .Z(n16007) );
  XOR U15842 ( .A(n15838), .B(n16010), .Z(n15831) );
  IV U15843 ( .A(n15837), .Z(n16010) );
  XNOR U15844 ( .A(n15834), .B(n16011), .Z(n15837) );
  XOR U15845 ( .A(n16012), .B(n16013), .Z(n15834) );
  ANDN U15846 ( .A(n16014), .B(n16015), .Z(n16013) );
  XNOR U15847 ( .A(n16012), .B(n16016), .Z(n16014) );
  XOR U15848 ( .A(n15845), .B(n16017), .Z(n15838) );
  IV U15849 ( .A(n15844), .Z(n16017) );
  XNOR U15850 ( .A(n15841), .B(n16018), .Z(n15844) );
  XOR U15851 ( .A(n16019), .B(n16020), .Z(n15841) );
  ANDN U15852 ( .A(n16021), .B(n16022), .Z(n16020) );
  XNOR U15853 ( .A(n16019), .B(n16023), .Z(n16021) );
  XOR U15854 ( .A(n15852), .B(n16024), .Z(n15845) );
  IV U15855 ( .A(n15851), .Z(n16024) );
  XNOR U15856 ( .A(n15848), .B(n16025), .Z(n15851) );
  XOR U15857 ( .A(n16026), .B(n16027), .Z(n15848) );
  ANDN U15858 ( .A(n16028), .B(n16029), .Z(n16027) );
  XNOR U15859 ( .A(n16026), .B(n16030), .Z(n16028) );
  XOR U15860 ( .A(n15859), .B(n16031), .Z(n15852) );
  IV U15861 ( .A(n15858), .Z(n16031) );
  XNOR U15862 ( .A(n15855), .B(n16032), .Z(n15858) );
  XOR U15863 ( .A(n16033), .B(n16034), .Z(n15855) );
  ANDN U15864 ( .A(n16035), .B(n16036), .Z(n16034) );
  XNOR U15865 ( .A(n16033), .B(n16037), .Z(n16035) );
  XOR U15866 ( .A(n15866), .B(n16038), .Z(n15859) );
  IV U15867 ( .A(n15865), .Z(n16038) );
  XNOR U15868 ( .A(n15862), .B(n16039), .Z(n15865) );
  XOR U15869 ( .A(n16040), .B(n16041), .Z(n15862) );
  ANDN U15870 ( .A(n16042), .B(n16043), .Z(n16041) );
  XNOR U15871 ( .A(n16040), .B(n16044), .Z(n16042) );
  XOR U15872 ( .A(n15873), .B(n16045), .Z(n15866) );
  IV U15873 ( .A(n15872), .Z(n16045) );
  XNOR U15874 ( .A(n15869), .B(n16046), .Z(n15872) );
  XOR U15875 ( .A(n16047), .B(n16048), .Z(n15869) );
  ANDN U15876 ( .A(n16049), .B(n16050), .Z(n16048) );
  XNOR U15877 ( .A(n16047), .B(n16051), .Z(n16049) );
  XOR U15878 ( .A(n15880), .B(n16052), .Z(n15873) );
  IV U15879 ( .A(n15879), .Z(n16052) );
  XNOR U15880 ( .A(n15876), .B(n16053), .Z(n15879) );
  XOR U15881 ( .A(n16054), .B(n16055), .Z(n15876) );
  ANDN U15882 ( .A(n16056), .B(n16057), .Z(n16055) );
  XNOR U15883 ( .A(n16054), .B(n16058), .Z(n16056) );
  XOR U15884 ( .A(n15887), .B(n16059), .Z(n15880) );
  IV U15885 ( .A(n15886), .Z(n16059) );
  XNOR U15886 ( .A(n15883), .B(n16060), .Z(n15886) );
  XOR U15887 ( .A(n16061), .B(n16062), .Z(n15883) );
  ANDN U15888 ( .A(n16063), .B(n16064), .Z(n16062) );
  XNOR U15889 ( .A(n16061), .B(n16065), .Z(n16063) );
  XOR U15890 ( .A(n15894), .B(n16066), .Z(n15887) );
  IV U15891 ( .A(n15893), .Z(n16066) );
  XNOR U15892 ( .A(n15890), .B(n16067), .Z(n15893) );
  XOR U15893 ( .A(n16068), .B(n16069), .Z(n15890) );
  ANDN U15894 ( .A(n16070), .B(n16071), .Z(n16069) );
  XNOR U15895 ( .A(n16068), .B(n16072), .Z(n16070) );
  XOR U15896 ( .A(n15901), .B(n16073), .Z(n15894) );
  IV U15897 ( .A(n15900), .Z(n16073) );
  XNOR U15898 ( .A(n15897), .B(n16074), .Z(n15900) );
  XOR U15899 ( .A(n16075), .B(n16076), .Z(n15897) );
  ANDN U15900 ( .A(n16077), .B(n16078), .Z(n16076) );
  XNOR U15901 ( .A(n16075), .B(n16079), .Z(n16077) );
  XOR U15902 ( .A(n15907), .B(n16080), .Z(n15901) );
  IV U15903 ( .A(n15906), .Z(n16080) );
  XNOR U15904 ( .A(n15903), .B(n16074), .Z(n15906) );
  AND U15905 ( .A(n16265), .B(n15896), .Z(n16074) );
  XOR U15906 ( .A(n16081), .B(n16082), .Z(n15903) );
  ANDN U15907 ( .A(n16083), .B(n16084), .Z(n16082) );
  XNOR U15908 ( .A(n16081), .B(n16085), .Z(n16083) );
  XOR U15909 ( .A(n15913), .B(n16086), .Z(n15907) );
  IV U15910 ( .A(n15912), .Z(n16086) );
  XNOR U15911 ( .A(n15909), .B(n16067), .Z(n15912) );
  AND U15912 ( .A(n16657), .B(n15553), .Z(n16067) );
  XOR U15913 ( .A(n16087), .B(n16088), .Z(n15909) );
  ANDN U15914 ( .A(n16089), .B(n16090), .Z(n16088) );
  XNOR U15915 ( .A(n16087), .B(n16091), .Z(n16089) );
  XOR U15916 ( .A(n15919), .B(n16092), .Z(n15913) );
  IV U15917 ( .A(n15918), .Z(n16092) );
  XNOR U15918 ( .A(n15915), .B(n16060), .Z(n15918) );
  AND U15919 ( .A(n17567), .B(n15236), .Z(n16060) );
  XOR U15920 ( .A(n16093), .B(n16094), .Z(n15915) );
  ANDN U15921 ( .A(n16095), .B(n16096), .Z(n16094) );
  XNOR U15922 ( .A(n16093), .B(n16097), .Z(n16095) );
  XOR U15923 ( .A(n15925), .B(n16098), .Z(n15919) );
  IV U15924 ( .A(n15924), .Z(n16098) );
  XNOR U15925 ( .A(n15921), .B(n16053), .Z(n15924) );
  AND U15926 ( .A(n17688), .B(n14945), .Z(n16053) );
  XOR U15927 ( .A(n16099), .B(n16100), .Z(n15921) );
  ANDN U15928 ( .A(n16101), .B(n16102), .Z(n16100) );
  XNOR U15929 ( .A(n16099), .B(n16103), .Z(n16101) );
  XOR U15930 ( .A(n15931), .B(n16104), .Z(n15925) );
  IV U15931 ( .A(n15930), .Z(n16104) );
  XNOR U15932 ( .A(n15927), .B(n16046), .Z(n15930) );
  AND U15933 ( .A(n17814), .B(n14680), .Z(n16046) );
  XOR U15934 ( .A(n16105), .B(n16106), .Z(n15927) );
  ANDN U15935 ( .A(n16107), .B(n16108), .Z(n16106) );
  XNOR U15936 ( .A(n16105), .B(n16109), .Z(n16107) );
  XOR U15937 ( .A(n15937), .B(n16110), .Z(n15931) );
  IV U15938 ( .A(n15936), .Z(n16110) );
  XNOR U15939 ( .A(n15933), .B(n16039), .Z(n15936) );
  AND U15940 ( .A(n17945), .B(n14441), .Z(n16039) );
  XOR U15941 ( .A(n16111), .B(n16112), .Z(n15933) );
  ANDN U15942 ( .A(n16113), .B(n16114), .Z(n16112) );
  XNOR U15943 ( .A(n16111), .B(n16115), .Z(n16113) );
  XOR U15944 ( .A(n15943), .B(n16116), .Z(n15937) );
  IV U15945 ( .A(n15942), .Z(n16116) );
  XNOR U15946 ( .A(n15939), .B(n16032), .Z(n15942) );
  AND U15947 ( .A(n18081), .B(n14228), .Z(n16032) );
  XOR U15948 ( .A(n16117), .B(n16118), .Z(n15939) );
  ANDN U15949 ( .A(n16119), .B(n16120), .Z(n16118) );
  XNOR U15950 ( .A(n16117), .B(n16121), .Z(n16119) );
  XOR U15951 ( .A(n15949), .B(n16122), .Z(n15943) );
  IV U15952 ( .A(n15948), .Z(n16122) );
  XNOR U15953 ( .A(n15945), .B(n16025), .Z(n15948) );
  AND U15954 ( .A(n18222), .B(n14041), .Z(n16025) );
  XOR U15955 ( .A(n16123), .B(n16124), .Z(n15945) );
  ANDN U15956 ( .A(n16125), .B(n16126), .Z(n16124) );
  XNOR U15957 ( .A(n16123), .B(n16127), .Z(n16125) );
  XOR U15958 ( .A(n15955), .B(n16128), .Z(n15949) );
  IV U15959 ( .A(n15954), .Z(n16128) );
  XNOR U15960 ( .A(n15951), .B(n16018), .Z(n15954) );
  AND U15961 ( .A(n18368), .B(n13880), .Z(n16018) );
  XOR U15962 ( .A(n16129), .B(n16130), .Z(n15951) );
  ANDN U15963 ( .A(n16131), .B(n16132), .Z(n16130) );
  XNOR U15964 ( .A(n16129), .B(n16133), .Z(n16131) );
  XOR U15965 ( .A(n15961), .B(n16134), .Z(n15955) );
  IV U15966 ( .A(n15960), .Z(n16134) );
  XNOR U15967 ( .A(n15957), .B(n16011), .Z(n15960) );
  AND U15968 ( .A(n18519), .B(n13745), .Z(n16011) );
  XOR U15969 ( .A(n16135), .B(n16136), .Z(n15957) );
  ANDN U15970 ( .A(n16137), .B(n16138), .Z(n16136) );
  XNOR U15971 ( .A(n16135), .B(n16139), .Z(n16137) );
  XOR U15972 ( .A(n15967), .B(n16140), .Z(n15961) );
  IV U15973 ( .A(n15966), .Z(n16140) );
  XNOR U15974 ( .A(n15963), .B(n16004), .Z(n15966) );
  AND U15975 ( .A(n18675), .B(n13636), .Z(n16004) );
  XOR U15976 ( .A(n16141), .B(n16142), .Z(n15963) );
  ANDN U15977 ( .A(n16143), .B(n16144), .Z(n16142) );
  XNOR U15978 ( .A(n16141), .B(n16145), .Z(n16143) );
  XOR U15979 ( .A(n15973), .B(n16146), .Z(n15967) );
  IV U15980 ( .A(n15972), .Z(n16146) );
  XNOR U15981 ( .A(n15969), .B(n15997), .Z(n15972) );
  AND U15982 ( .A(n18836), .B(n13553), .Z(n15997) );
  XOR U15983 ( .A(n16147), .B(n16148), .Z(n15969) );
  ANDN U15984 ( .A(n16149), .B(n16150), .Z(n16148) );
  XNOR U15985 ( .A(n16147), .B(n16151), .Z(n16149) );
  XOR U15986 ( .A(n15979), .B(n16152), .Z(n15973) );
  IV U15987 ( .A(n15978), .Z(n16152) );
  XNOR U15988 ( .A(n15975), .B(n15990), .Z(n15978) );
  AND U15989 ( .A(n19002), .B(n13496), .Z(n15990) );
  XOR U15990 ( .A(n16153), .B(n16154), .Z(n15975) );
  ANDN U15991 ( .A(n16155), .B(n16156), .Z(n16154) );
  XNOR U15992 ( .A(n16153), .B(n16157), .Z(n16155) );
  XOR U15993 ( .A(n15984), .B(n16158), .Z(n15979) );
  IV U15994 ( .A(n15983), .Z(n16158) );
  XNOR U15995 ( .A(n15980), .B(n15988), .Z(n15983) );
  AND U15996 ( .A(n13470), .B(n19173), .Z(n15988) );
  XOR U15997 ( .A(n16159), .B(n16160), .Z(n15980) );
  ANDN U15998 ( .A(n16161), .B(n16162), .Z(n16160) );
  XNOR U15999 ( .A(n16159), .B(n16163), .Z(n16161) );
  XNOR U16000 ( .A(n16164), .B(n16165), .Z(n15984) );
  ANDN U16001 ( .A(n16166), .B(n16167), .Z(n16165) );
  XNOR U16002 ( .A(n16164), .B(n16168), .Z(n16166) );
  XOR U16003 ( .A(n16169), .B(n16170), .Z(n15985) );
  ANDN U16004 ( .A(n16171), .B(n8864), .Z(n16170) );
  XNOR U16005 ( .A(n16169), .B(n16172), .Z(n8864) );
  XNOR U16006 ( .A(n16169), .B(n8862), .Z(n16171) );
  XOR U16007 ( .A(n15995), .B(n16173), .Z(n8862) );
  IV U16008 ( .A(n15994), .Z(n16173) );
  XNOR U16009 ( .A(n15991), .B(n16174), .Z(n15994) );
  XOR U16010 ( .A(n16175), .B(n16176), .Z(n15991) );
  ANDN U16011 ( .A(n16177), .B(n16178), .Z(n16176) );
  XNOR U16012 ( .A(n16175), .B(n16179), .Z(n16177) );
  XOR U16013 ( .A(n16002), .B(n16180), .Z(n15995) );
  IV U16014 ( .A(n16001), .Z(n16180) );
  XNOR U16015 ( .A(n15998), .B(n16181), .Z(n16001) );
  XOR U16016 ( .A(n16182), .B(n16183), .Z(n15998) );
  ANDN U16017 ( .A(n16184), .B(n16185), .Z(n16183) );
  XNOR U16018 ( .A(n16182), .B(n16186), .Z(n16184) );
  XOR U16019 ( .A(n16009), .B(n16187), .Z(n16002) );
  IV U16020 ( .A(n16008), .Z(n16187) );
  XNOR U16021 ( .A(n16005), .B(n16188), .Z(n16008) );
  XOR U16022 ( .A(n16189), .B(n16190), .Z(n16005) );
  ANDN U16023 ( .A(n16191), .B(n16192), .Z(n16190) );
  XNOR U16024 ( .A(n16189), .B(n16193), .Z(n16191) );
  XOR U16025 ( .A(n16016), .B(n16194), .Z(n16009) );
  IV U16026 ( .A(n16015), .Z(n16194) );
  XNOR U16027 ( .A(n16012), .B(n16195), .Z(n16015) );
  XOR U16028 ( .A(n16196), .B(n16197), .Z(n16012) );
  ANDN U16029 ( .A(n16198), .B(n16199), .Z(n16197) );
  XNOR U16030 ( .A(n16196), .B(n16200), .Z(n16198) );
  XOR U16031 ( .A(n16023), .B(n16201), .Z(n16016) );
  IV U16032 ( .A(n16022), .Z(n16201) );
  XNOR U16033 ( .A(n16019), .B(n16202), .Z(n16022) );
  XOR U16034 ( .A(n16203), .B(n16204), .Z(n16019) );
  ANDN U16035 ( .A(n16205), .B(n16206), .Z(n16204) );
  XNOR U16036 ( .A(n16203), .B(n16207), .Z(n16205) );
  XOR U16037 ( .A(n16030), .B(n16208), .Z(n16023) );
  IV U16038 ( .A(n16029), .Z(n16208) );
  XNOR U16039 ( .A(n16026), .B(n16209), .Z(n16029) );
  XOR U16040 ( .A(n16210), .B(n16211), .Z(n16026) );
  ANDN U16041 ( .A(n16212), .B(n16213), .Z(n16211) );
  XNOR U16042 ( .A(n16210), .B(n16214), .Z(n16212) );
  XOR U16043 ( .A(n16037), .B(n16215), .Z(n16030) );
  IV U16044 ( .A(n16036), .Z(n16215) );
  XNOR U16045 ( .A(n16033), .B(n16216), .Z(n16036) );
  XOR U16046 ( .A(n16217), .B(n16218), .Z(n16033) );
  ANDN U16047 ( .A(n16219), .B(n16220), .Z(n16218) );
  XNOR U16048 ( .A(n16217), .B(n16221), .Z(n16219) );
  XOR U16049 ( .A(n16044), .B(n16222), .Z(n16037) );
  IV U16050 ( .A(n16043), .Z(n16222) );
  XNOR U16051 ( .A(n16040), .B(n16223), .Z(n16043) );
  XOR U16052 ( .A(n16224), .B(n16225), .Z(n16040) );
  ANDN U16053 ( .A(n16226), .B(n16227), .Z(n16225) );
  XNOR U16054 ( .A(n16224), .B(n16228), .Z(n16226) );
  XOR U16055 ( .A(n16051), .B(n16229), .Z(n16044) );
  IV U16056 ( .A(n16050), .Z(n16229) );
  XNOR U16057 ( .A(n16047), .B(n16230), .Z(n16050) );
  XOR U16058 ( .A(n16231), .B(n16232), .Z(n16047) );
  ANDN U16059 ( .A(n16233), .B(n16234), .Z(n16232) );
  XNOR U16060 ( .A(n16231), .B(n16235), .Z(n16233) );
  XOR U16061 ( .A(n16058), .B(n16236), .Z(n16051) );
  IV U16062 ( .A(n16057), .Z(n16236) );
  XNOR U16063 ( .A(n16054), .B(n16237), .Z(n16057) );
  XOR U16064 ( .A(n16238), .B(n16239), .Z(n16054) );
  ANDN U16065 ( .A(n16240), .B(n16241), .Z(n16239) );
  XNOR U16066 ( .A(n16238), .B(n16242), .Z(n16240) );
  XOR U16067 ( .A(n16065), .B(n16243), .Z(n16058) );
  IV U16068 ( .A(n16064), .Z(n16243) );
  XNOR U16069 ( .A(n16061), .B(n16244), .Z(n16064) );
  XOR U16070 ( .A(n16245), .B(n16246), .Z(n16061) );
  ANDN U16071 ( .A(n16247), .B(n16248), .Z(n16246) );
  XNOR U16072 ( .A(n16245), .B(n16249), .Z(n16247) );
  XOR U16073 ( .A(n16072), .B(n16250), .Z(n16065) );
  IV U16074 ( .A(n16071), .Z(n16250) );
  XNOR U16075 ( .A(n16068), .B(n16251), .Z(n16071) );
  XOR U16076 ( .A(n16252), .B(n16253), .Z(n16068) );
  ANDN U16077 ( .A(n16254), .B(n16255), .Z(n16253) );
  XNOR U16078 ( .A(n16252), .B(n16256), .Z(n16254) );
  XOR U16079 ( .A(n16079), .B(n16257), .Z(n16072) );
  IV U16080 ( .A(n16078), .Z(n16257) );
  XNOR U16081 ( .A(n16075), .B(n16258), .Z(n16078) );
  XOR U16082 ( .A(n16259), .B(n16260), .Z(n16075) );
  ANDN U16083 ( .A(n16261), .B(n16262), .Z(n16260) );
  XNOR U16084 ( .A(n16259), .B(n16263), .Z(n16261) );
  XOR U16085 ( .A(n16085), .B(n16264), .Z(n16079) );
  IV U16086 ( .A(n16084), .Z(n16264) );
  XNOR U16087 ( .A(n16081), .B(n16265), .Z(n16084) );
  XOR U16088 ( .A(n16266), .B(n16267), .Z(n16081) );
  ANDN U16089 ( .A(n16268), .B(n16269), .Z(n16267) );
  XNOR U16090 ( .A(n16266), .B(n16270), .Z(n16268) );
  XOR U16091 ( .A(n16091), .B(n16271), .Z(n16085) );
  IV U16092 ( .A(n16090), .Z(n16271) );
  XNOR U16093 ( .A(n16087), .B(n16258), .Z(n16090) );
  AND U16094 ( .A(n16657), .B(n15896), .Z(n16258) );
  XOR U16095 ( .A(n16272), .B(n16273), .Z(n16087) );
  ANDN U16096 ( .A(n16274), .B(n16275), .Z(n16273) );
  XNOR U16097 ( .A(n16272), .B(n16276), .Z(n16274) );
  XOR U16098 ( .A(n16097), .B(n16277), .Z(n16091) );
  IV U16099 ( .A(n16096), .Z(n16277) );
  XNOR U16100 ( .A(n16093), .B(n16251), .Z(n16096) );
  AND U16101 ( .A(n17567), .B(n15553), .Z(n16251) );
  XOR U16102 ( .A(n16278), .B(n16279), .Z(n16093) );
  ANDN U16103 ( .A(n16280), .B(n16281), .Z(n16279) );
  XNOR U16104 ( .A(n16278), .B(n16282), .Z(n16280) );
  XOR U16105 ( .A(n16103), .B(n16283), .Z(n16097) );
  IV U16106 ( .A(n16102), .Z(n16283) );
  XNOR U16107 ( .A(n16099), .B(n16244), .Z(n16102) );
  AND U16108 ( .A(n17688), .B(n15236), .Z(n16244) );
  XOR U16109 ( .A(n16284), .B(n16285), .Z(n16099) );
  ANDN U16110 ( .A(n16286), .B(n16287), .Z(n16285) );
  XNOR U16111 ( .A(n16284), .B(n16288), .Z(n16286) );
  XOR U16112 ( .A(n16109), .B(n16289), .Z(n16103) );
  IV U16113 ( .A(n16108), .Z(n16289) );
  XNOR U16114 ( .A(n16105), .B(n16237), .Z(n16108) );
  AND U16115 ( .A(n17814), .B(n14945), .Z(n16237) );
  XOR U16116 ( .A(n16290), .B(n16291), .Z(n16105) );
  ANDN U16117 ( .A(n16292), .B(n16293), .Z(n16291) );
  XNOR U16118 ( .A(n16290), .B(n16294), .Z(n16292) );
  XOR U16119 ( .A(n16115), .B(n16295), .Z(n16109) );
  IV U16120 ( .A(n16114), .Z(n16295) );
  XNOR U16121 ( .A(n16111), .B(n16230), .Z(n16114) );
  AND U16122 ( .A(n17945), .B(n14680), .Z(n16230) );
  XOR U16123 ( .A(n16296), .B(n16297), .Z(n16111) );
  ANDN U16124 ( .A(n16298), .B(n16299), .Z(n16297) );
  XNOR U16125 ( .A(n16296), .B(n16300), .Z(n16298) );
  XOR U16126 ( .A(n16121), .B(n16301), .Z(n16115) );
  IV U16127 ( .A(n16120), .Z(n16301) );
  XNOR U16128 ( .A(n16117), .B(n16223), .Z(n16120) );
  AND U16129 ( .A(n18081), .B(n14441), .Z(n16223) );
  XOR U16130 ( .A(n16302), .B(n16303), .Z(n16117) );
  ANDN U16131 ( .A(n16304), .B(n16305), .Z(n16303) );
  XNOR U16132 ( .A(n16302), .B(n16306), .Z(n16304) );
  XOR U16133 ( .A(n16127), .B(n16307), .Z(n16121) );
  IV U16134 ( .A(n16126), .Z(n16307) );
  XNOR U16135 ( .A(n16123), .B(n16216), .Z(n16126) );
  AND U16136 ( .A(n18222), .B(n14228), .Z(n16216) );
  XOR U16137 ( .A(n16308), .B(n16309), .Z(n16123) );
  ANDN U16138 ( .A(n16310), .B(n16311), .Z(n16309) );
  XNOR U16139 ( .A(n16308), .B(n16312), .Z(n16310) );
  XOR U16140 ( .A(n16133), .B(n16313), .Z(n16127) );
  IV U16141 ( .A(n16132), .Z(n16313) );
  XNOR U16142 ( .A(n16129), .B(n16209), .Z(n16132) );
  AND U16143 ( .A(n18368), .B(n14041), .Z(n16209) );
  XOR U16144 ( .A(n16314), .B(n16315), .Z(n16129) );
  ANDN U16145 ( .A(n16316), .B(n16317), .Z(n16315) );
  XNOR U16146 ( .A(n16314), .B(n16318), .Z(n16316) );
  XOR U16147 ( .A(n16139), .B(n16319), .Z(n16133) );
  IV U16148 ( .A(n16138), .Z(n16319) );
  XNOR U16149 ( .A(n16135), .B(n16202), .Z(n16138) );
  AND U16150 ( .A(n18519), .B(n13880), .Z(n16202) );
  XOR U16151 ( .A(n16320), .B(n16321), .Z(n16135) );
  ANDN U16152 ( .A(n16322), .B(n16323), .Z(n16321) );
  XNOR U16153 ( .A(n16320), .B(n16324), .Z(n16322) );
  XOR U16154 ( .A(n16145), .B(n16325), .Z(n16139) );
  IV U16155 ( .A(n16144), .Z(n16325) );
  XNOR U16156 ( .A(n16141), .B(n16195), .Z(n16144) );
  AND U16157 ( .A(n18675), .B(n13745), .Z(n16195) );
  XOR U16158 ( .A(n16326), .B(n16327), .Z(n16141) );
  ANDN U16159 ( .A(n16328), .B(n16329), .Z(n16327) );
  XNOR U16160 ( .A(n16326), .B(n16330), .Z(n16328) );
  XOR U16161 ( .A(n16151), .B(n16331), .Z(n16145) );
  IV U16162 ( .A(n16150), .Z(n16331) );
  XNOR U16163 ( .A(n16147), .B(n16188), .Z(n16150) );
  AND U16164 ( .A(n18836), .B(n13636), .Z(n16188) );
  XOR U16165 ( .A(n16332), .B(n16333), .Z(n16147) );
  ANDN U16166 ( .A(n16334), .B(n16335), .Z(n16333) );
  XNOR U16167 ( .A(n16332), .B(n16336), .Z(n16334) );
  XOR U16168 ( .A(n16157), .B(n16337), .Z(n16151) );
  IV U16169 ( .A(n16156), .Z(n16337) );
  XNOR U16170 ( .A(n16153), .B(n16181), .Z(n16156) );
  AND U16171 ( .A(n19002), .B(n13553), .Z(n16181) );
  XOR U16172 ( .A(n16338), .B(n16339), .Z(n16153) );
  ANDN U16173 ( .A(n16340), .B(n16341), .Z(n16339) );
  XNOR U16174 ( .A(n16338), .B(n16342), .Z(n16340) );
  XOR U16175 ( .A(n16163), .B(n16343), .Z(n16157) );
  IV U16176 ( .A(n16162), .Z(n16343) );
  XNOR U16177 ( .A(n16159), .B(n16174), .Z(n16162) );
  AND U16178 ( .A(n19173), .B(n13496), .Z(n16174) );
  XOR U16179 ( .A(n16344), .B(n16345), .Z(n16159) );
  ANDN U16180 ( .A(n16346), .B(n16347), .Z(n16345) );
  XNOR U16181 ( .A(n16344), .B(n16348), .Z(n16346) );
  XOR U16182 ( .A(n16168), .B(n16349), .Z(n16163) );
  IV U16183 ( .A(n16167), .Z(n16349) );
  XNOR U16184 ( .A(n16164), .B(n16172), .Z(n16167) );
  AND U16185 ( .A(n13470), .B(n19349), .Z(n16172) );
  XOR U16186 ( .A(n16350), .B(n16351), .Z(n16164) );
  ANDN U16187 ( .A(n16352), .B(n16353), .Z(n16351) );
  XNOR U16188 ( .A(n16350), .B(n16354), .Z(n16352) );
  XNOR U16189 ( .A(n16355), .B(n16356), .Z(n16168) );
  ANDN U16190 ( .A(n16357), .B(n16358), .Z(n16356) );
  XNOR U16191 ( .A(n16355), .B(n16359), .Z(n16357) );
  XOR U16192 ( .A(n16360), .B(n16361), .Z(n16169) );
  ANDN U16193 ( .A(n16362), .B(n9089), .Z(n16361) );
  XNOR U16194 ( .A(n16360), .B(n16363), .Z(n9089) );
  XNOR U16195 ( .A(n16360), .B(n9087), .Z(n16362) );
  XOR U16196 ( .A(n16179), .B(n16364), .Z(n9087) );
  IV U16197 ( .A(n16178), .Z(n16364) );
  XNOR U16198 ( .A(n16175), .B(n16365), .Z(n16178) );
  XOR U16199 ( .A(n16366), .B(n16367), .Z(n16175) );
  ANDN U16200 ( .A(n16368), .B(n16369), .Z(n16367) );
  XNOR U16201 ( .A(n16366), .B(n16370), .Z(n16368) );
  XOR U16202 ( .A(n16186), .B(n16371), .Z(n16179) );
  IV U16203 ( .A(n16185), .Z(n16371) );
  XNOR U16204 ( .A(n16182), .B(n16372), .Z(n16185) );
  XOR U16205 ( .A(n16373), .B(n16374), .Z(n16182) );
  ANDN U16206 ( .A(n16375), .B(n16376), .Z(n16374) );
  XNOR U16207 ( .A(n16373), .B(n16377), .Z(n16375) );
  XOR U16208 ( .A(n16193), .B(n16378), .Z(n16186) );
  IV U16209 ( .A(n16192), .Z(n16378) );
  XNOR U16210 ( .A(n16189), .B(n16379), .Z(n16192) );
  XOR U16211 ( .A(n16380), .B(n16381), .Z(n16189) );
  ANDN U16212 ( .A(n16382), .B(n16383), .Z(n16381) );
  XNOR U16213 ( .A(n16380), .B(n16384), .Z(n16382) );
  XOR U16214 ( .A(n16200), .B(n16385), .Z(n16193) );
  IV U16215 ( .A(n16199), .Z(n16385) );
  XNOR U16216 ( .A(n16196), .B(n16386), .Z(n16199) );
  XOR U16217 ( .A(n16387), .B(n16388), .Z(n16196) );
  ANDN U16218 ( .A(n16389), .B(n16390), .Z(n16388) );
  XNOR U16219 ( .A(n16387), .B(n16391), .Z(n16389) );
  XOR U16220 ( .A(n16207), .B(n16392), .Z(n16200) );
  IV U16221 ( .A(n16206), .Z(n16392) );
  XNOR U16222 ( .A(n16203), .B(n16393), .Z(n16206) );
  XOR U16223 ( .A(n16394), .B(n16395), .Z(n16203) );
  ANDN U16224 ( .A(n16396), .B(n16397), .Z(n16395) );
  XNOR U16225 ( .A(n16394), .B(n16398), .Z(n16396) );
  XOR U16226 ( .A(n16214), .B(n16399), .Z(n16207) );
  IV U16227 ( .A(n16213), .Z(n16399) );
  XNOR U16228 ( .A(n16210), .B(n16400), .Z(n16213) );
  XOR U16229 ( .A(n16401), .B(n16402), .Z(n16210) );
  ANDN U16230 ( .A(n16403), .B(n16404), .Z(n16402) );
  XNOR U16231 ( .A(n16401), .B(n16405), .Z(n16403) );
  XOR U16232 ( .A(n16221), .B(n16406), .Z(n16214) );
  IV U16233 ( .A(n16220), .Z(n16406) );
  XNOR U16234 ( .A(n16217), .B(n16407), .Z(n16220) );
  XOR U16235 ( .A(n16408), .B(n16409), .Z(n16217) );
  ANDN U16236 ( .A(n16410), .B(n16411), .Z(n16409) );
  XNOR U16237 ( .A(n16408), .B(n16412), .Z(n16410) );
  XOR U16238 ( .A(n16228), .B(n16413), .Z(n16221) );
  IV U16239 ( .A(n16227), .Z(n16413) );
  XNOR U16240 ( .A(n16224), .B(n16414), .Z(n16227) );
  XOR U16241 ( .A(n16415), .B(n16416), .Z(n16224) );
  ANDN U16242 ( .A(n16417), .B(n16418), .Z(n16416) );
  XNOR U16243 ( .A(n16415), .B(n16419), .Z(n16417) );
  XOR U16244 ( .A(n16235), .B(n16420), .Z(n16228) );
  IV U16245 ( .A(n16234), .Z(n16420) );
  XNOR U16246 ( .A(n16231), .B(n16421), .Z(n16234) );
  XOR U16247 ( .A(n16422), .B(n16423), .Z(n16231) );
  ANDN U16248 ( .A(n16424), .B(n16425), .Z(n16423) );
  XNOR U16249 ( .A(n16422), .B(n16426), .Z(n16424) );
  XOR U16250 ( .A(n16242), .B(n16427), .Z(n16235) );
  IV U16251 ( .A(n16241), .Z(n16427) );
  XNOR U16252 ( .A(n16238), .B(n16428), .Z(n16241) );
  XOR U16253 ( .A(n16429), .B(n16430), .Z(n16238) );
  ANDN U16254 ( .A(n16431), .B(n16432), .Z(n16430) );
  XNOR U16255 ( .A(n16429), .B(n16433), .Z(n16431) );
  XOR U16256 ( .A(n16249), .B(n16434), .Z(n16242) );
  IV U16257 ( .A(n16248), .Z(n16434) );
  XNOR U16258 ( .A(n16245), .B(n16435), .Z(n16248) );
  XOR U16259 ( .A(n16436), .B(n16437), .Z(n16245) );
  ANDN U16260 ( .A(n16438), .B(n16439), .Z(n16437) );
  XNOR U16261 ( .A(n16436), .B(n16440), .Z(n16438) );
  XOR U16262 ( .A(n16256), .B(n16441), .Z(n16249) );
  IV U16263 ( .A(n16255), .Z(n16441) );
  XNOR U16264 ( .A(n16252), .B(n16442), .Z(n16255) );
  XOR U16265 ( .A(n16443), .B(n16444), .Z(n16252) );
  ANDN U16266 ( .A(n16445), .B(n16446), .Z(n16444) );
  XNOR U16267 ( .A(n16443), .B(n16447), .Z(n16445) );
  XOR U16268 ( .A(n16263), .B(n16448), .Z(n16256) );
  IV U16269 ( .A(n16262), .Z(n16448) );
  XNOR U16270 ( .A(n16259), .B(n16449), .Z(n16262) );
  XOR U16271 ( .A(n16450), .B(n16451), .Z(n16259) );
  ANDN U16272 ( .A(n16452), .B(n16453), .Z(n16451) );
  XNOR U16273 ( .A(n16450), .B(n16454), .Z(n16452) );
  XOR U16274 ( .A(n16270), .B(n16455), .Z(n16263) );
  IV U16275 ( .A(n16269), .Z(n16455) );
  XNOR U16276 ( .A(n16266), .B(n16456), .Z(n16269) );
  XOR U16277 ( .A(n16457), .B(n16458), .Z(n16266) );
  ANDN U16278 ( .A(n16459), .B(n16460), .Z(n16458) );
  XNOR U16279 ( .A(n16457), .B(n16461), .Z(n16459) );
  XOR U16280 ( .A(n16276), .B(n16462), .Z(n16270) );
  IV U16281 ( .A(n16275), .Z(n16462) );
  XNOR U16282 ( .A(n16272), .B(n16456), .Z(n16275) );
  AND U16283 ( .A(n16657), .B(n16265), .Z(n16456) );
  XOR U16284 ( .A(n16463), .B(n16464), .Z(n16272) );
  ANDN U16285 ( .A(n16465), .B(n16466), .Z(n16464) );
  XNOR U16286 ( .A(n16463), .B(n16467), .Z(n16465) );
  XOR U16287 ( .A(n16282), .B(n16468), .Z(n16276) );
  IV U16288 ( .A(n16281), .Z(n16468) );
  XNOR U16289 ( .A(n16278), .B(n16449), .Z(n16281) );
  AND U16290 ( .A(n17567), .B(n15896), .Z(n16449) );
  XOR U16291 ( .A(n16469), .B(n16470), .Z(n16278) );
  ANDN U16292 ( .A(n16471), .B(n16472), .Z(n16470) );
  XNOR U16293 ( .A(n16469), .B(n16473), .Z(n16471) );
  XOR U16294 ( .A(n16288), .B(n16474), .Z(n16282) );
  IV U16295 ( .A(n16287), .Z(n16474) );
  XNOR U16296 ( .A(n16284), .B(n16442), .Z(n16287) );
  AND U16297 ( .A(n17688), .B(n15553), .Z(n16442) );
  XOR U16298 ( .A(n16475), .B(n16476), .Z(n16284) );
  ANDN U16299 ( .A(n16477), .B(n16478), .Z(n16476) );
  XNOR U16300 ( .A(n16475), .B(n16479), .Z(n16477) );
  XOR U16301 ( .A(n16294), .B(n16480), .Z(n16288) );
  IV U16302 ( .A(n16293), .Z(n16480) );
  XNOR U16303 ( .A(n16290), .B(n16435), .Z(n16293) );
  AND U16304 ( .A(n17814), .B(n15236), .Z(n16435) );
  XOR U16305 ( .A(n16481), .B(n16482), .Z(n16290) );
  ANDN U16306 ( .A(n16483), .B(n16484), .Z(n16482) );
  XNOR U16307 ( .A(n16481), .B(n16485), .Z(n16483) );
  XOR U16308 ( .A(n16300), .B(n16486), .Z(n16294) );
  IV U16309 ( .A(n16299), .Z(n16486) );
  XNOR U16310 ( .A(n16296), .B(n16428), .Z(n16299) );
  AND U16311 ( .A(n17945), .B(n14945), .Z(n16428) );
  XOR U16312 ( .A(n16487), .B(n16488), .Z(n16296) );
  ANDN U16313 ( .A(n16489), .B(n16490), .Z(n16488) );
  XNOR U16314 ( .A(n16487), .B(n16491), .Z(n16489) );
  XOR U16315 ( .A(n16306), .B(n16492), .Z(n16300) );
  IV U16316 ( .A(n16305), .Z(n16492) );
  XNOR U16317 ( .A(n16302), .B(n16421), .Z(n16305) );
  AND U16318 ( .A(n18081), .B(n14680), .Z(n16421) );
  XOR U16319 ( .A(n16493), .B(n16494), .Z(n16302) );
  ANDN U16320 ( .A(n16495), .B(n16496), .Z(n16494) );
  XNOR U16321 ( .A(n16493), .B(n16497), .Z(n16495) );
  XOR U16322 ( .A(n16312), .B(n16498), .Z(n16306) );
  IV U16323 ( .A(n16311), .Z(n16498) );
  XNOR U16324 ( .A(n16308), .B(n16414), .Z(n16311) );
  AND U16325 ( .A(n18222), .B(n14441), .Z(n16414) );
  XOR U16326 ( .A(n16499), .B(n16500), .Z(n16308) );
  ANDN U16327 ( .A(n16501), .B(n16502), .Z(n16500) );
  XNOR U16328 ( .A(n16499), .B(n16503), .Z(n16501) );
  XOR U16329 ( .A(n16318), .B(n16504), .Z(n16312) );
  IV U16330 ( .A(n16317), .Z(n16504) );
  XNOR U16331 ( .A(n16314), .B(n16407), .Z(n16317) );
  AND U16332 ( .A(n18368), .B(n14228), .Z(n16407) );
  XOR U16333 ( .A(n16505), .B(n16506), .Z(n16314) );
  ANDN U16334 ( .A(n16507), .B(n16508), .Z(n16506) );
  XNOR U16335 ( .A(n16505), .B(n16509), .Z(n16507) );
  XOR U16336 ( .A(n16324), .B(n16510), .Z(n16318) );
  IV U16337 ( .A(n16323), .Z(n16510) );
  XNOR U16338 ( .A(n16320), .B(n16400), .Z(n16323) );
  AND U16339 ( .A(n18519), .B(n14041), .Z(n16400) );
  XOR U16340 ( .A(n16511), .B(n16512), .Z(n16320) );
  ANDN U16341 ( .A(n16513), .B(n16514), .Z(n16512) );
  XNOR U16342 ( .A(n16511), .B(n16515), .Z(n16513) );
  XOR U16343 ( .A(n16330), .B(n16516), .Z(n16324) );
  IV U16344 ( .A(n16329), .Z(n16516) );
  XNOR U16345 ( .A(n16326), .B(n16393), .Z(n16329) );
  AND U16346 ( .A(n18675), .B(n13880), .Z(n16393) );
  XOR U16347 ( .A(n16517), .B(n16518), .Z(n16326) );
  ANDN U16348 ( .A(n16519), .B(n16520), .Z(n16518) );
  XNOR U16349 ( .A(n16517), .B(n16521), .Z(n16519) );
  XOR U16350 ( .A(n16336), .B(n16522), .Z(n16330) );
  IV U16351 ( .A(n16335), .Z(n16522) );
  XNOR U16352 ( .A(n16332), .B(n16386), .Z(n16335) );
  AND U16353 ( .A(n18836), .B(n13745), .Z(n16386) );
  XOR U16354 ( .A(n16523), .B(n16524), .Z(n16332) );
  ANDN U16355 ( .A(n16525), .B(n16526), .Z(n16524) );
  XNOR U16356 ( .A(n16523), .B(n16527), .Z(n16525) );
  XOR U16357 ( .A(n16342), .B(n16528), .Z(n16336) );
  IV U16358 ( .A(n16341), .Z(n16528) );
  XNOR U16359 ( .A(n16338), .B(n16379), .Z(n16341) );
  AND U16360 ( .A(n19002), .B(n13636), .Z(n16379) );
  XOR U16361 ( .A(n16529), .B(n16530), .Z(n16338) );
  ANDN U16362 ( .A(n16531), .B(n16532), .Z(n16530) );
  XNOR U16363 ( .A(n16529), .B(n16533), .Z(n16531) );
  XOR U16364 ( .A(n16348), .B(n16534), .Z(n16342) );
  IV U16365 ( .A(n16347), .Z(n16534) );
  XNOR U16366 ( .A(n16344), .B(n16372), .Z(n16347) );
  AND U16367 ( .A(n19173), .B(n13553), .Z(n16372) );
  XOR U16368 ( .A(n16535), .B(n16536), .Z(n16344) );
  ANDN U16369 ( .A(n16537), .B(n16538), .Z(n16536) );
  XNOR U16370 ( .A(n16535), .B(n16539), .Z(n16537) );
  XOR U16371 ( .A(n16354), .B(n16540), .Z(n16348) );
  IV U16372 ( .A(n16353), .Z(n16540) );
  XNOR U16373 ( .A(n16350), .B(n16365), .Z(n16353) );
  AND U16374 ( .A(n19349), .B(n13496), .Z(n16365) );
  XOR U16375 ( .A(n16541), .B(n16542), .Z(n16350) );
  ANDN U16376 ( .A(n16543), .B(n16544), .Z(n16542) );
  XNOR U16377 ( .A(n16541), .B(n16545), .Z(n16543) );
  XOR U16378 ( .A(n16359), .B(n16546), .Z(n16354) );
  IV U16379 ( .A(n16358), .Z(n16546) );
  XNOR U16380 ( .A(n16355), .B(n16363), .Z(n16358) );
  AND U16381 ( .A(n13470), .B(n19478), .Z(n16363) );
  XOR U16382 ( .A(n16547), .B(n16548), .Z(n16355) );
  ANDN U16383 ( .A(n16549), .B(n16550), .Z(n16548) );
  XOR U16384 ( .A(n16547), .B(n16551), .Z(n16549) );
  XNOR U16385 ( .A(n16552), .B(n16553), .Z(n16359) );
  ANDN U16386 ( .A(n16552), .B(n16554), .Z(n16553) );
  XOR U16387 ( .A(n16555), .B(n16556), .Z(n16360) );
  NANDN U16388 ( .B(n9308), .A(n16557), .Z(n16555) );
  XOR U16389 ( .A(n16556), .B(n9306), .Z(n16557) );
  XOR U16390 ( .A(n16370), .B(n16558), .Z(n9306) );
  IV U16391 ( .A(n16369), .Z(n16558) );
  XNOR U16392 ( .A(n16366), .B(n16559), .Z(n16369) );
  XOR U16393 ( .A(n16560), .B(n16561), .Z(n16366) );
  NANDN U16394 ( .B(n16562), .A(n16563), .Z(n16560) );
  XOR U16395 ( .A(n16561), .B(n16564), .Z(n16563) );
  XOR U16396 ( .A(n16377), .B(n16565), .Z(n16370) );
  IV U16397 ( .A(n16376), .Z(n16565) );
  XNOR U16398 ( .A(n16373), .B(n16566), .Z(n16376) );
  XOR U16399 ( .A(n16567), .B(n16568), .Z(n16373) );
  ANDN U16400 ( .A(n16569), .B(n16570), .Z(n16568) );
  XNOR U16401 ( .A(n16567), .B(n16571), .Z(n16569) );
  XOR U16402 ( .A(n16384), .B(n16572), .Z(n16377) );
  IV U16403 ( .A(n16383), .Z(n16572) );
  XNOR U16404 ( .A(n16380), .B(n16573), .Z(n16383) );
  XOR U16405 ( .A(n16574), .B(n16575), .Z(n16380) );
  ANDN U16406 ( .A(n16576), .B(n16577), .Z(n16575) );
  XNOR U16407 ( .A(n16574), .B(n16578), .Z(n16576) );
  XOR U16408 ( .A(n16391), .B(n16579), .Z(n16384) );
  IV U16409 ( .A(n16390), .Z(n16579) );
  XNOR U16410 ( .A(n16387), .B(n16580), .Z(n16390) );
  XOR U16411 ( .A(n16581), .B(n16582), .Z(n16387) );
  ANDN U16412 ( .A(n16583), .B(n16584), .Z(n16582) );
  XNOR U16413 ( .A(n16581), .B(n16585), .Z(n16583) );
  XOR U16414 ( .A(n16398), .B(n16586), .Z(n16391) );
  IV U16415 ( .A(n16397), .Z(n16586) );
  XNOR U16416 ( .A(n16394), .B(n16587), .Z(n16397) );
  XOR U16417 ( .A(n16588), .B(n16589), .Z(n16394) );
  ANDN U16418 ( .A(n16590), .B(n16591), .Z(n16589) );
  XNOR U16419 ( .A(n16588), .B(n16592), .Z(n16590) );
  XOR U16420 ( .A(n16405), .B(n16593), .Z(n16398) );
  IV U16421 ( .A(n16404), .Z(n16593) );
  XNOR U16422 ( .A(n16401), .B(n16594), .Z(n16404) );
  XOR U16423 ( .A(n16595), .B(n16596), .Z(n16401) );
  ANDN U16424 ( .A(n16597), .B(n16598), .Z(n16596) );
  XNOR U16425 ( .A(n16595), .B(n16599), .Z(n16597) );
  XOR U16426 ( .A(n16412), .B(n16600), .Z(n16405) );
  IV U16427 ( .A(n16411), .Z(n16600) );
  XNOR U16428 ( .A(n16408), .B(n16601), .Z(n16411) );
  XOR U16429 ( .A(n16602), .B(n16603), .Z(n16408) );
  ANDN U16430 ( .A(n16604), .B(n16605), .Z(n16603) );
  XNOR U16431 ( .A(n16602), .B(n16606), .Z(n16604) );
  XOR U16432 ( .A(n16419), .B(n16607), .Z(n16412) );
  IV U16433 ( .A(n16418), .Z(n16607) );
  XNOR U16434 ( .A(n16415), .B(n16608), .Z(n16418) );
  XOR U16435 ( .A(n16609), .B(n16610), .Z(n16415) );
  ANDN U16436 ( .A(n16611), .B(n16612), .Z(n16610) );
  XNOR U16437 ( .A(n16609), .B(n16613), .Z(n16611) );
  XOR U16438 ( .A(n16426), .B(n16614), .Z(n16419) );
  IV U16439 ( .A(n16425), .Z(n16614) );
  XNOR U16440 ( .A(n16422), .B(n16615), .Z(n16425) );
  XOR U16441 ( .A(n16616), .B(n16617), .Z(n16422) );
  ANDN U16442 ( .A(n16618), .B(n16619), .Z(n16617) );
  XNOR U16443 ( .A(n16616), .B(n16620), .Z(n16618) );
  XOR U16444 ( .A(n16433), .B(n16621), .Z(n16426) );
  IV U16445 ( .A(n16432), .Z(n16621) );
  XNOR U16446 ( .A(n16429), .B(n16622), .Z(n16432) );
  XOR U16447 ( .A(n16623), .B(n16624), .Z(n16429) );
  ANDN U16448 ( .A(n16625), .B(n16626), .Z(n16624) );
  XNOR U16449 ( .A(n16623), .B(n16627), .Z(n16625) );
  XOR U16450 ( .A(n16440), .B(n16628), .Z(n16433) );
  IV U16451 ( .A(n16439), .Z(n16628) );
  XNOR U16452 ( .A(n16436), .B(n16629), .Z(n16439) );
  XOR U16453 ( .A(n16630), .B(n16631), .Z(n16436) );
  ANDN U16454 ( .A(n16632), .B(n16633), .Z(n16631) );
  XNOR U16455 ( .A(n16630), .B(n16634), .Z(n16632) );
  XOR U16456 ( .A(n16447), .B(n16635), .Z(n16440) );
  IV U16457 ( .A(n16446), .Z(n16635) );
  XNOR U16458 ( .A(n16443), .B(n16636), .Z(n16446) );
  XOR U16459 ( .A(n16637), .B(n16638), .Z(n16443) );
  ANDN U16460 ( .A(n16639), .B(n16640), .Z(n16638) );
  XNOR U16461 ( .A(n16637), .B(n16641), .Z(n16639) );
  XOR U16462 ( .A(n16454), .B(n16642), .Z(n16447) );
  IV U16463 ( .A(n16453), .Z(n16642) );
  XNOR U16464 ( .A(n16450), .B(n16643), .Z(n16453) );
  XOR U16465 ( .A(n16644), .B(n16645), .Z(n16450) );
  ANDN U16466 ( .A(n16646), .B(n16647), .Z(n16645) );
  XNOR U16467 ( .A(n16644), .B(n16648), .Z(n16646) );
  XOR U16468 ( .A(n16461), .B(n16649), .Z(n16454) );
  IV U16469 ( .A(n16460), .Z(n16649) );
  XNOR U16470 ( .A(n16457), .B(n16650), .Z(n16460) );
  XOR U16471 ( .A(n16651), .B(n16652), .Z(n16457) );
  ANDN U16472 ( .A(n16653), .B(n16654), .Z(n16652) );
  XNOR U16473 ( .A(n16651), .B(n16655), .Z(n16653) );
  XOR U16474 ( .A(n16467), .B(n16656), .Z(n16461) );
  IV U16475 ( .A(n16466), .Z(n16656) );
  XNOR U16476 ( .A(n16463), .B(n16657), .Z(n16466) );
  XOR U16477 ( .A(n16658), .B(n16659), .Z(n16463) );
  ANDN U16478 ( .A(n16660), .B(n16661), .Z(n16659) );
  XNOR U16479 ( .A(n16658), .B(n16662), .Z(n16660) );
  XOR U16480 ( .A(n16473), .B(n16663), .Z(n16467) );
  IV U16481 ( .A(n16472), .Z(n16663) );
  XNOR U16482 ( .A(n16469), .B(n16650), .Z(n16472) );
  AND U16483 ( .A(n17567), .B(n16265), .Z(n16650) );
  XOR U16484 ( .A(n16664), .B(n16665), .Z(n16469) );
  ANDN U16485 ( .A(n16666), .B(n16667), .Z(n16665) );
  XNOR U16486 ( .A(n16664), .B(n16668), .Z(n16666) );
  XOR U16487 ( .A(n16479), .B(n16669), .Z(n16473) );
  IV U16488 ( .A(n16478), .Z(n16669) );
  XNOR U16489 ( .A(n16475), .B(n16643), .Z(n16478) );
  AND U16490 ( .A(n17688), .B(n15896), .Z(n16643) );
  XOR U16491 ( .A(n16670), .B(n16671), .Z(n16475) );
  ANDN U16492 ( .A(n16672), .B(n16673), .Z(n16671) );
  XNOR U16493 ( .A(n16670), .B(n16674), .Z(n16672) );
  XOR U16494 ( .A(n16485), .B(n16675), .Z(n16479) );
  IV U16495 ( .A(n16484), .Z(n16675) );
  XNOR U16496 ( .A(n16481), .B(n16636), .Z(n16484) );
  AND U16497 ( .A(n17814), .B(n15553), .Z(n16636) );
  XOR U16498 ( .A(n16676), .B(n16677), .Z(n16481) );
  ANDN U16499 ( .A(n16678), .B(n16679), .Z(n16677) );
  XNOR U16500 ( .A(n16676), .B(n16680), .Z(n16678) );
  XOR U16501 ( .A(n16491), .B(n16681), .Z(n16485) );
  IV U16502 ( .A(n16490), .Z(n16681) );
  XNOR U16503 ( .A(n16487), .B(n16629), .Z(n16490) );
  AND U16504 ( .A(n17945), .B(n15236), .Z(n16629) );
  XOR U16505 ( .A(n16682), .B(n16683), .Z(n16487) );
  ANDN U16506 ( .A(n16684), .B(n16685), .Z(n16683) );
  XNOR U16507 ( .A(n16682), .B(n16686), .Z(n16684) );
  XOR U16508 ( .A(n16497), .B(n16687), .Z(n16491) );
  IV U16509 ( .A(n16496), .Z(n16687) );
  XNOR U16510 ( .A(n16493), .B(n16622), .Z(n16496) );
  AND U16511 ( .A(n18081), .B(n14945), .Z(n16622) );
  XOR U16512 ( .A(n16688), .B(n16689), .Z(n16493) );
  ANDN U16513 ( .A(n16690), .B(n16691), .Z(n16689) );
  XNOR U16514 ( .A(n16688), .B(n16692), .Z(n16690) );
  XOR U16515 ( .A(n16503), .B(n16693), .Z(n16497) );
  IV U16516 ( .A(n16502), .Z(n16693) );
  XNOR U16517 ( .A(n16499), .B(n16615), .Z(n16502) );
  AND U16518 ( .A(n18222), .B(n14680), .Z(n16615) );
  XOR U16519 ( .A(n16694), .B(n16695), .Z(n16499) );
  ANDN U16520 ( .A(n16696), .B(n16697), .Z(n16695) );
  XNOR U16521 ( .A(n16694), .B(n16698), .Z(n16696) );
  XOR U16522 ( .A(n16509), .B(n16699), .Z(n16503) );
  IV U16523 ( .A(n16508), .Z(n16699) );
  XNOR U16524 ( .A(n16505), .B(n16608), .Z(n16508) );
  AND U16525 ( .A(n18368), .B(n14441), .Z(n16608) );
  XOR U16526 ( .A(n16700), .B(n16701), .Z(n16505) );
  ANDN U16527 ( .A(n16702), .B(n16703), .Z(n16701) );
  XNOR U16528 ( .A(n16700), .B(n16704), .Z(n16702) );
  XOR U16529 ( .A(n16515), .B(n16705), .Z(n16509) );
  IV U16530 ( .A(n16514), .Z(n16705) );
  XNOR U16531 ( .A(n16511), .B(n16601), .Z(n16514) );
  AND U16532 ( .A(n18519), .B(n14228), .Z(n16601) );
  XOR U16533 ( .A(n16706), .B(n16707), .Z(n16511) );
  ANDN U16534 ( .A(n16708), .B(n16709), .Z(n16707) );
  XNOR U16535 ( .A(n16706), .B(n16710), .Z(n16708) );
  XOR U16536 ( .A(n16521), .B(n16711), .Z(n16515) );
  IV U16537 ( .A(n16520), .Z(n16711) );
  XNOR U16538 ( .A(n16517), .B(n16594), .Z(n16520) );
  AND U16539 ( .A(n18675), .B(n14041), .Z(n16594) );
  XOR U16540 ( .A(n16712), .B(n16713), .Z(n16517) );
  ANDN U16541 ( .A(n16714), .B(n16715), .Z(n16713) );
  XNOR U16542 ( .A(n16712), .B(n16716), .Z(n16714) );
  XOR U16543 ( .A(n16527), .B(n16717), .Z(n16521) );
  IV U16544 ( .A(n16526), .Z(n16717) );
  XNOR U16545 ( .A(n16523), .B(n16587), .Z(n16526) );
  AND U16546 ( .A(n18836), .B(n13880), .Z(n16587) );
  XOR U16547 ( .A(n16718), .B(n16719), .Z(n16523) );
  ANDN U16548 ( .A(n16720), .B(n16721), .Z(n16719) );
  XNOR U16549 ( .A(n16718), .B(n16722), .Z(n16720) );
  XOR U16550 ( .A(n16533), .B(n16723), .Z(n16527) );
  IV U16551 ( .A(n16532), .Z(n16723) );
  XNOR U16552 ( .A(n16529), .B(n16580), .Z(n16532) );
  AND U16553 ( .A(n19002), .B(n13745), .Z(n16580) );
  XOR U16554 ( .A(n16724), .B(n16725), .Z(n16529) );
  ANDN U16555 ( .A(n16726), .B(n16727), .Z(n16725) );
  XNOR U16556 ( .A(n16724), .B(n16728), .Z(n16726) );
  XOR U16557 ( .A(n16539), .B(n16729), .Z(n16533) );
  IV U16558 ( .A(n16538), .Z(n16729) );
  XNOR U16559 ( .A(n16535), .B(n16573), .Z(n16538) );
  AND U16560 ( .A(n19173), .B(n13636), .Z(n16573) );
  XOR U16561 ( .A(n16730), .B(n16731), .Z(n16535) );
  ANDN U16562 ( .A(n16732), .B(n16733), .Z(n16731) );
  XNOR U16563 ( .A(n16730), .B(n16734), .Z(n16732) );
  XOR U16564 ( .A(n16545), .B(n16735), .Z(n16539) );
  IV U16565 ( .A(n16544), .Z(n16735) );
  XNOR U16566 ( .A(n16541), .B(n16566), .Z(n16544) );
  AND U16567 ( .A(n19349), .B(n13553), .Z(n16566) );
  XOR U16568 ( .A(n16736), .B(n16737), .Z(n16541) );
  ANDN U16569 ( .A(n16738), .B(n16739), .Z(n16737) );
  XNOR U16570 ( .A(n16736), .B(n16740), .Z(n16738) );
  XOR U16571 ( .A(n16551), .B(n16550), .Z(n16545) );
  XNOR U16572 ( .A(n16547), .B(n16559), .Z(n16550) );
  AND U16573 ( .A(n19478), .B(n13496), .Z(n16559) );
  XOR U16574 ( .A(n16741), .B(n16742), .Z(n16547) );
  ANDN U16575 ( .A(n16743), .B(n16744), .Z(n16742) );
  XNOR U16576 ( .A(n16741), .B(n16745), .Z(n16743) );
  IV U16577 ( .A(n16554), .Z(n16551) );
  XNOR U16578 ( .A(n16552), .B(n16746), .Z(n16554) );
  AND U16579 ( .A(n13470), .B(n16747), .Z(n16746) );
  XOR U16580 ( .A(n16748), .B(n16749), .Z(n16552) );
  ANDN U16581 ( .A(n16750), .B(n16751), .Z(n16749) );
  XNOR U16582 ( .A(n9519), .B(n16748), .Z(n16750) );
  XNOR U16583 ( .A(n16752), .B(n16556), .Z(n9308) );
  OR U16584 ( .A(n9518), .B(n9519), .Z(n16556) );
  XOR U16585 ( .A(n16564), .B(n16753), .Z(n9518) );
  IV U16586 ( .A(n16562), .Z(n16753) );
  XNOR U16587 ( .A(n16754), .B(n16561), .Z(n16562) );
  OR U16588 ( .A(n9723), .B(n9724), .Z(n16561) );
  XOR U16589 ( .A(n16755), .B(n16756), .Z(n9723) );
  IV U16590 ( .A(n16757), .Z(n16756) );
  NAND U16591 ( .A(n16747), .B(n13496), .Z(n16754) );
  XOR U16592 ( .A(n16571), .B(n16758), .Z(n16564) );
  IV U16593 ( .A(n16570), .Z(n16758) );
  XNOR U16594 ( .A(n16567), .B(n16759), .Z(n16570) );
  XOR U16595 ( .A(n16760), .B(n16761), .Z(n16567) );
  NANDN U16596 ( .B(n16757), .A(n16762), .Z(n16760) );
  XOR U16597 ( .A(n16761), .B(n16755), .Z(n16762) );
  XOR U16598 ( .A(n16763), .B(n16764), .Z(n16755) );
  IV U16599 ( .A(n16765), .Z(n16764) );
  XNOR U16600 ( .A(n16766), .B(n16761), .Z(n16757) );
  OR U16601 ( .A(n9921), .B(n9922), .Z(n16761) );
  XOR U16602 ( .A(n16767), .B(n16768), .Z(n9921) );
  IV U16603 ( .A(n16769), .Z(n16768) );
  NAND U16604 ( .A(n16747), .B(n13553), .Z(n16766) );
  XOR U16605 ( .A(n16578), .B(n16770), .Z(n16571) );
  IV U16606 ( .A(n16577), .Z(n16770) );
  XNOR U16607 ( .A(n16574), .B(n16771), .Z(n16577) );
  XOR U16608 ( .A(n16772), .B(n16773), .Z(n16574) );
  ANDN U16609 ( .A(n16774), .B(n16765), .Z(n16773) );
  XNOR U16610 ( .A(n16772), .B(n16775), .Z(n16765) );
  XNOR U16611 ( .A(n16772), .B(n16763), .Z(n16774) );
  XOR U16612 ( .A(n16776), .B(n16777), .Z(n16763) );
  IV U16613 ( .A(n16778), .Z(n16777) );
  XOR U16614 ( .A(n16779), .B(n16780), .Z(n16772) );
  NANDN U16615 ( .B(n16769), .A(n16781), .Z(n16779) );
  XOR U16616 ( .A(n16780), .B(n16767), .Z(n16781) );
  XOR U16617 ( .A(n16782), .B(n16783), .Z(n16767) );
  IV U16618 ( .A(n16784), .Z(n16783) );
  XNOR U16619 ( .A(n16785), .B(n16780), .Z(n16769) );
  OR U16620 ( .A(n10113), .B(n10114), .Z(n16780) );
  XOR U16621 ( .A(n16786), .B(n16787), .Z(n10113) );
  IV U16622 ( .A(n16788), .Z(n16787) );
  NAND U16623 ( .A(n16747), .B(n13636), .Z(n16785) );
  XOR U16624 ( .A(n16585), .B(n16789), .Z(n16578) );
  IV U16625 ( .A(n16584), .Z(n16789) );
  XNOR U16626 ( .A(n16581), .B(n16790), .Z(n16584) );
  XOR U16627 ( .A(n16791), .B(n16792), .Z(n16581) );
  ANDN U16628 ( .A(n16793), .B(n16778), .Z(n16792) );
  XNOR U16629 ( .A(n16791), .B(n16794), .Z(n16778) );
  XNOR U16630 ( .A(n16791), .B(n16776), .Z(n16793) );
  XOR U16631 ( .A(n16795), .B(n16796), .Z(n16776) );
  IV U16632 ( .A(n16797), .Z(n16796) );
  XOR U16633 ( .A(n16798), .B(n16799), .Z(n16791) );
  ANDN U16634 ( .A(n16800), .B(n16784), .Z(n16799) );
  XNOR U16635 ( .A(n16798), .B(n16801), .Z(n16784) );
  XNOR U16636 ( .A(n16798), .B(n16782), .Z(n16800) );
  XOR U16637 ( .A(n16802), .B(n16803), .Z(n16782) );
  IV U16638 ( .A(n16804), .Z(n16803) );
  XOR U16639 ( .A(n16805), .B(n16806), .Z(n16798) );
  NANDN U16640 ( .B(n16788), .A(n16807), .Z(n16805) );
  XOR U16641 ( .A(n16806), .B(n16786), .Z(n16807) );
  XOR U16642 ( .A(n16808), .B(n16809), .Z(n16786) );
  IV U16643 ( .A(n16810), .Z(n16809) );
  XNOR U16644 ( .A(n16811), .B(n16806), .Z(n16788) );
  OR U16645 ( .A(n10298), .B(n10299), .Z(n16806) );
  XOR U16646 ( .A(n16812), .B(n16813), .Z(n10298) );
  IV U16647 ( .A(n16814), .Z(n16813) );
  NAND U16648 ( .A(n16747), .B(n13745), .Z(n16811) );
  XOR U16649 ( .A(n16592), .B(n16815), .Z(n16585) );
  IV U16650 ( .A(n16591), .Z(n16815) );
  XNOR U16651 ( .A(n16588), .B(n16816), .Z(n16591) );
  XOR U16652 ( .A(n16817), .B(n16818), .Z(n16588) );
  ANDN U16653 ( .A(n16819), .B(n16797), .Z(n16818) );
  XNOR U16654 ( .A(n16817), .B(n16820), .Z(n16797) );
  XNOR U16655 ( .A(n16817), .B(n16795), .Z(n16819) );
  XOR U16656 ( .A(n16821), .B(n16822), .Z(n16795) );
  IV U16657 ( .A(n16823), .Z(n16822) );
  XOR U16658 ( .A(n16824), .B(n16825), .Z(n16817) );
  ANDN U16659 ( .A(n16826), .B(n16804), .Z(n16825) );
  XNOR U16660 ( .A(n16824), .B(n16827), .Z(n16804) );
  XNOR U16661 ( .A(n16824), .B(n16802), .Z(n16826) );
  XOR U16662 ( .A(n16828), .B(n16829), .Z(n16802) );
  IV U16663 ( .A(n16830), .Z(n16829) );
  XOR U16664 ( .A(n16831), .B(n16832), .Z(n16824) );
  ANDN U16665 ( .A(n16833), .B(n16810), .Z(n16832) );
  XNOR U16666 ( .A(n16831), .B(n16834), .Z(n16810) );
  XNOR U16667 ( .A(n16831), .B(n16808), .Z(n16833) );
  XOR U16668 ( .A(n16835), .B(n16836), .Z(n16808) );
  IV U16669 ( .A(n16837), .Z(n16836) );
  XOR U16670 ( .A(n16838), .B(n16839), .Z(n16831) );
  NANDN U16671 ( .B(n16814), .A(n16840), .Z(n16838) );
  XOR U16672 ( .A(n16839), .B(n16812), .Z(n16840) );
  XOR U16673 ( .A(n16841), .B(n16842), .Z(n16812) );
  IV U16674 ( .A(n16843), .Z(n16842) );
  XNOR U16675 ( .A(n16844), .B(n16839), .Z(n16814) );
  OR U16676 ( .A(n10477), .B(n10478), .Z(n16839) );
  XOR U16677 ( .A(n16845), .B(n16846), .Z(n10477) );
  IV U16678 ( .A(n16847), .Z(n16846) );
  NAND U16679 ( .A(n16747), .B(n13880), .Z(n16844) );
  XOR U16680 ( .A(n16599), .B(n16848), .Z(n16592) );
  IV U16681 ( .A(n16598), .Z(n16848) );
  XNOR U16682 ( .A(n16595), .B(n16849), .Z(n16598) );
  XOR U16683 ( .A(n16850), .B(n16851), .Z(n16595) );
  ANDN U16684 ( .A(n16852), .B(n16823), .Z(n16851) );
  XNOR U16685 ( .A(n16850), .B(n16853), .Z(n16823) );
  XNOR U16686 ( .A(n16850), .B(n16821), .Z(n16852) );
  XOR U16687 ( .A(n16854), .B(n16855), .Z(n16821) );
  IV U16688 ( .A(n16856), .Z(n16855) );
  XOR U16689 ( .A(n16857), .B(n16858), .Z(n16850) );
  ANDN U16690 ( .A(n16859), .B(n16830), .Z(n16858) );
  XNOR U16691 ( .A(n16857), .B(n16860), .Z(n16830) );
  XNOR U16692 ( .A(n16857), .B(n16828), .Z(n16859) );
  XOR U16693 ( .A(n16861), .B(n16862), .Z(n16828) );
  IV U16694 ( .A(n16863), .Z(n16862) );
  XOR U16695 ( .A(n16864), .B(n16865), .Z(n16857) );
  ANDN U16696 ( .A(n16866), .B(n16837), .Z(n16865) );
  XNOR U16697 ( .A(n16864), .B(n16867), .Z(n16837) );
  XNOR U16698 ( .A(n16864), .B(n16835), .Z(n16866) );
  XOR U16699 ( .A(n16868), .B(n16869), .Z(n16835) );
  IV U16700 ( .A(n16870), .Z(n16869) );
  XOR U16701 ( .A(n16871), .B(n16872), .Z(n16864) );
  ANDN U16702 ( .A(n16873), .B(n16843), .Z(n16872) );
  XNOR U16703 ( .A(n16871), .B(n16874), .Z(n16843) );
  XNOR U16704 ( .A(n16871), .B(n16841), .Z(n16873) );
  XOR U16705 ( .A(n16875), .B(n16876), .Z(n16841) );
  IV U16706 ( .A(n16877), .Z(n16876) );
  XOR U16707 ( .A(n16878), .B(n16879), .Z(n16871) );
  NANDN U16708 ( .B(n16847), .A(n16880), .Z(n16878) );
  XOR U16709 ( .A(n16879), .B(n16845), .Z(n16880) );
  XOR U16710 ( .A(n16881), .B(n16882), .Z(n16845) );
  IV U16711 ( .A(n16883), .Z(n16882) );
  XNOR U16712 ( .A(n16884), .B(n16879), .Z(n16847) );
  OR U16713 ( .A(n10649), .B(n10650), .Z(n16879) );
  XOR U16714 ( .A(n16885), .B(n16886), .Z(n10649) );
  IV U16715 ( .A(n16887), .Z(n16886) );
  NAND U16716 ( .A(n16747), .B(n14041), .Z(n16884) );
  XOR U16717 ( .A(n16606), .B(n16888), .Z(n16599) );
  IV U16718 ( .A(n16605), .Z(n16888) );
  XNOR U16719 ( .A(n16602), .B(n16889), .Z(n16605) );
  XOR U16720 ( .A(n16890), .B(n16891), .Z(n16602) );
  ANDN U16721 ( .A(n16892), .B(n16856), .Z(n16891) );
  XNOR U16722 ( .A(n16890), .B(n16893), .Z(n16856) );
  XNOR U16723 ( .A(n16890), .B(n16854), .Z(n16892) );
  XOR U16724 ( .A(n16894), .B(n16895), .Z(n16854) );
  IV U16725 ( .A(n16896), .Z(n16895) );
  XOR U16726 ( .A(n16897), .B(n16898), .Z(n16890) );
  ANDN U16727 ( .A(n16899), .B(n16863), .Z(n16898) );
  XNOR U16728 ( .A(n16897), .B(n16900), .Z(n16863) );
  XNOR U16729 ( .A(n16897), .B(n16861), .Z(n16899) );
  XOR U16730 ( .A(n16901), .B(n16902), .Z(n16861) );
  IV U16731 ( .A(n16903), .Z(n16902) );
  XOR U16732 ( .A(n16904), .B(n16905), .Z(n16897) );
  ANDN U16733 ( .A(n16906), .B(n16870), .Z(n16905) );
  XNOR U16734 ( .A(n16904), .B(n16907), .Z(n16870) );
  XNOR U16735 ( .A(n16904), .B(n16868), .Z(n16906) );
  XOR U16736 ( .A(n16908), .B(n16909), .Z(n16868) );
  IV U16737 ( .A(n16910), .Z(n16909) );
  XOR U16738 ( .A(n16911), .B(n16912), .Z(n16904) );
  ANDN U16739 ( .A(n16913), .B(n16877), .Z(n16912) );
  XNOR U16740 ( .A(n16911), .B(n16914), .Z(n16877) );
  XNOR U16741 ( .A(n16911), .B(n16875), .Z(n16913) );
  XOR U16742 ( .A(n16915), .B(n16916), .Z(n16875) );
  IV U16743 ( .A(n16917), .Z(n16916) );
  XOR U16744 ( .A(n16918), .B(n16919), .Z(n16911) );
  ANDN U16745 ( .A(n16920), .B(n16883), .Z(n16919) );
  XNOR U16746 ( .A(n16918), .B(n16921), .Z(n16883) );
  XNOR U16747 ( .A(n16918), .B(n16881), .Z(n16920) );
  XOR U16748 ( .A(n16922), .B(n16923), .Z(n16881) );
  IV U16749 ( .A(n16924), .Z(n16923) );
  XOR U16750 ( .A(n16925), .B(n16926), .Z(n16918) );
  NANDN U16751 ( .B(n16887), .A(n16927), .Z(n16925) );
  XOR U16752 ( .A(n16926), .B(n16885), .Z(n16927) );
  XOR U16753 ( .A(n16928), .B(n16929), .Z(n16885) );
  IV U16754 ( .A(n16930), .Z(n16929) );
  XNOR U16755 ( .A(n16931), .B(n16926), .Z(n16887) );
  OR U16756 ( .A(n10815), .B(n10816), .Z(n16926) );
  XOR U16757 ( .A(n16932), .B(n16933), .Z(n10815) );
  IV U16758 ( .A(n16934), .Z(n16933) );
  NAND U16759 ( .A(n16747), .B(n14228), .Z(n16931) );
  XOR U16760 ( .A(n16613), .B(n16935), .Z(n16606) );
  IV U16761 ( .A(n16612), .Z(n16935) );
  XNOR U16762 ( .A(n16609), .B(n16936), .Z(n16612) );
  XOR U16763 ( .A(n16937), .B(n16938), .Z(n16609) );
  ANDN U16764 ( .A(n16939), .B(n16896), .Z(n16938) );
  XNOR U16765 ( .A(n16937), .B(n16940), .Z(n16896) );
  XNOR U16766 ( .A(n16937), .B(n16894), .Z(n16939) );
  XOR U16767 ( .A(n16941), .B(n16942), .Z(n16894) );
  IV U16768 ( .A(n16943), .Z(n16942) );
  XOR U16769 ( .A(n16944), .B(n16945), .Z(n16937) );
  ANDN U16770 ( .A(n16946), .B(n16903), .Z(n16945) );
  XNOR U16771 ( .A(n16944), .B(n16947), .Z(n16903) );
  XNOR U16772 ( .A(n16944), .B(n16901), .Z(n16946) );
  XOR U16773 ( .A(n16948), .B(n16949), .Z(n16901) );
  IV U16774 ( .A(n16950), .Z(n16949) );
  XOR U16775 ( .A(n16951), .B(n16952), .Z(n16944) );
  ANDN U16776 ( .A(n16953), .B(n16910), .Z(n16952) );
  XNOR U16777 ( .A(n16951), .B(n16954), .Z(n16910) );
  XNOR U16778 ( .A(n16951), .B(n16908), .Z(n16953) );
  XOR U16779 ( .A(n16955), .B(n16956), .Z(n16908) );
  IV U16780 ( .A(n16957), .Z(n16956) );
  XOR U16781 ( .A(n16958), .B(n16959), .Z(n16951) );
  ANDN U16782 ( .A(n16960), .B(n16917), .Z(n16959) );
  XNOR U16783 ( .A(n16958), .B(n16961), .Z(n16917) );
  XNOR U16784 ( .A(n16958), .B(n16915), .Z(n16960) );
  XOR U16785 ( .A(n16962), .B(n16963), .Z(n16915) );
  IV U16786 ( .A(n16964), .Z(n16963) );
  XOR U16787 ( .A(n16965), .B(n16966), .Z(n16958) );
  ANDN U16788 ( .A(n16967), .B(n16924), .Z(n16966) );
  XNOR U16789 ( .A(n16965), .B(n16968), .Z(n16924) );
  XNOR U16790 ( .A(n16965), .B(n16922), .Z(n16967) );
  XOR U16791 ( .A(n16969), .B(n16970), .Z(n16922) );
  IV U16792 ( .A(n16971), .Z(n16970) );
  XOR U16793 ( .A(n16972), .B(n16973), .Z(n16965) );
  ANDN U16794 ( .A(n16974), .B(n16930), .Z(n16973) );
  XNOR U16795 ( .A(n16972), .B(n16975), .Z(n16930) );
  XNOR U16796 ( .A(n16972), .B(n16928), .Z(n16974) );
  XOR U16797 ( .A(n16976), .B(n16977), .Z(n16928) );
  IV U16798 ( .A(n16978), .Z(n16977) );
  XOR U16799 ( .A(n16979), .B(n16980), .Z(n16972) );
  NANDN U16800 ( .B(n16934), .A(n16981), .Z(n16979) );
  XOR U16801 ( .A(n16980), .B(n16932), .Z(n16981) );
  XOR U16802 ( .A(n16982), .B(n16983), .Z(n16932) );
  IV U16803 ( .A(n16984), .Z(n16983) );
  XNOR U16804 ( .A(n16985), .B(n16980), .Z(n16934) );
  OR U16805 ( .A(n10974), .B(n10975), .Z(n16980) );
  XOR U16806 ( .A(n16986), .B(n16987), .Z(n10974) );
  IV U16807 ( .A(n16988), .Z(n16987) );
  NAND U16808 ( .A(n16747), .B(n14441), .Z(n16985) );
  XOR U16809 ( .A(n16620), .B(n16989), .Z(n16613) );
  IV U16810 ( .A(n16619), .Z(n16989) );
  XNOR U16811 ( .A(n16616), .B(n16990), .Z(n16619) );
  XOR U16812 ( .A(n16991), .B(n16992), .Z(n16616) );
  ANDN U16813 ( .A(n16993), .B(n16943), .Z(n16992) );
  XNOR U16814 ( .A(n16991), .B(n16994), .Z(n16943) );
  XNOR U16815 ( .A(n16991), .B(n16941), .Z(n16993) );
  XOR U16816 ( .A(n16995), .B(n16996), .Z(n16941) );
  IV U16817 ( .A(n16997), .Z(n16996) );
  XOR U16818 ( .A(n16998), .B(n16999), .Z(n16991) );
  ANDN U16819 ( .A(n17000), .B(n16950), .Z(n16999) );
  XNOR U16820 ( .A(n16998), .B(n17001), .Z(n16950) );
  XNOR U16821 ( .A(n16998), .B(n16948), .Z(n17000) );
  XOR U16822 ( .A(n17002), .B(n17003), .Z(n16948) );
  IV U16823 ( .A(n17004), .Z(n17003) );
  XOR U16824 ( .A(n17005), .B(n17006), .Z(n16998) );
  ANDN U16825 ( .A(n17007), .B(n16957), .Z(n17006) );
  XNOR U16826 ( .A(n17005), .B(n17008), .Z(n16957) );
  XNOR U16827 ( .A(n17005), .B(n16955), .Z(n17007) );
  XOR U16828 ( .A(n17009), .B(n17010), .Z(n16955) );
  IV U16829 ( .A(n17011), .Z(n17010) );
  XOR U16830 ( .A(n17012), .B(n17013), .Z(n17005) );
  ANDN U16831 ( .A(n17014), .B(n16964), .Z(n17013) );
  XNOR U16832 ( .A(n17012), .B(n17015), .Z(n16964) );
  XNOR U16833 ( .A(n17012), .B(n16962), .Z(n17014) );
  XOR U16834 ( .A(n17016), .B(n17017), .Z(n16962) );
  IV U16835 ( .A(n17018), .Z(n17017) );
  XOR U16836 ( .A(n17019), .B(n17020), .Z(n17012) );
  ANDN U16837 ( .A(n17021), .B(n16971), .Z(n17020) );
  XNOR U16838 ( .A(n17019), .B(n17022), .Z(n16971) );
  XNOR U16839 ( .A(n17019), .B(n16969), .Z(n17021) );
  XOR U16840 ( .A(n17023), .B(n17024), .Z(n16969) );
  IV U16841 ( .A(n17025), .Z(n17024) );
  XOR U16842 ( .A(n17026), .B(n17027), .Z(n17019) );
  ANDN U16843 ( .A(n17028), .B(n16978), .Z(n17027) );
  XNOR U16844 ( .A(n17026), .B(n17029), .Z(n16978) );
  XNOR U16845 ( .A(n17026), .B(n16976), .Z(n17028) );
  XOR U16846 ( .A(n17030), .B(n17031), .Z(n16976) );
  IV U16847 ( .A(n17032), .Z(n17031) );
  XOR U16848 ( .A(n17033), .B(n17034), .Z(n17026) );
  ANDN U16849 ( .A(n17035), .B(n16984), .Z(n17034) );
  XNOR U16850 ( .A(n17033), .B(n17036), .Z(n16984) );
  XNOR U16851 ( .A(n17033), .B(n16982), .Z(n17035) );
  XOR U16852 ( .A(n17037), .B(n17038), .Z(n16982) );
  IV U16853 ( .A(n17039), .Z(n17038) );
  XOR U16854 ( .A(n17040), .B(n17041), .Z(n17033) );
  NANDN U16855 ( .B(n16988), .A(n17042), .Z(n17040) );
  XOR U16856 ( .A(n17041), .B(n16986), .Z(n17042) );
  XOR U16857 ( .A(n17043), .B(n17044), .Z(n16986) );
  IV U16858 ( .A(n17045), .Z(n17044) );
  XNOR U16859 ( .A(n17046), .B(n17041), .Z(n16988) );
  OR U16860 ( .A(n11127), .B(n11128), .Z(n17041) );
  XOR U16861 ( .A(n17047), .B(n17048), .Z(n11127) );
  IV U16862 ( .A(n17049), .Z(n17048) );
  NAND U16863 ( .A(n16747), .B(n14680), .Z(n17046) );
  XOR U16864 ( .A(n16627), .B(n17050), .Z(n16620) );
  IV U16865 ( .A(n16626), .Z(n17050) );
  XNOR U16866 ( .A(n16623), .B(n17051), .Z(n16626) );
  XOR U16867 ( .A(n17052), .B(n17053), .Z(n16623) );
  ANDN U16868 ( .A(n17054), .B(n16997), .Z(n17053) );
  XNOR U16869 ( .A(n17052), .B(n17055), .Z(n16997) );
  XNOR U16870 ( .A(n17052), .B(n16995), .Z(n17054) );
  XOR U16871 ( .A(n17056), .B(n17057), .Z(n16995) );
  IV U16872 ( .A(n17058), .Z(n17057) );
  XOR U16873 ( .A(n17059), .B(n17060), .Z(n17052) );
  ANDN U16874 ( .A(n17061), .B(n17004), .Z(n17060) );
  XNOR U16875 ( .A(n17059), .B(n17062), .Z(n17004) );
  XNOR U16876 ( .A(n17059), .B(n17002), .Z(n17061) );
  XOR U16877 ( .A(n17063), .B(n17064), .Z(n17002) );
  IV U16878 ( .A(n17065), .Z(n17064) );
  XOR U16879 ( .A(n17066), .B(n17067), .Z(n17059) );
  ANDN U16880 ( .A(n17068), .B(n17011), .Z(n17067) );
  XNOR U16881 ( .A(n17066), .B(n17069), .Z(n17011) );
  XNOR U16882 ( .A(n17066), .B(n17009), .Z(n17068) );
  XOR U16883 ( .A(n17070), .B(n17071), .Z(n17009) );
  IV U16884 ( .A(n17072), .Z(n17071) );
  XOR U16885 ( .A(n17073), .B(n17074), .Z(n17066) );
  ANDN U16886 ( .A(n17075), .B(n17018), .Z(n17074) );
  XNOR U16887 ( .A(n17073), .B(n17076), .Z(n17018) );
  XNOR U16888 ( .A(n17073), .B(n17016), .Z(n17075) );
  XOR U16889 ( .A(n17077), .B(n17078), .Z(n17016) );
  IV U16890 ( .A(n17079), .Z(n17078) );
  XOR U16891 ( .A(n17080), .B(n17081), .Z(n17073) );
  ANDN U16892 ( .A(n17082), .B(n17025), .Z(n17081) );
  XNOR U16893 ( .A(n17080), .B(n17083), .Z(n17025) );
  XNOR U16894 ( .A(n17080), .B(n17023), .Z(n17082) );
  XOR U16895 ( .A(n17084), .B(n17085), .Z(n17023) );
  IV U16896 ( .A(n17086), .Z(n17085) );
  XOR U16897 ( .A(n17087), .B(n17088), .Z(n17080) );
  ANDN U16898 ( .A(n17089), .B(n17032), .Z(n17088) );
  XNOR U16899 ( .A(n17087), .B(n17090), .Z(n17032) );
  XNOR U16900 ( .A(n17087), .B(n17030), .Z(n17089) );
  XOR U16901 ( .A(n17091), .B(n17092), .Z(n17030) );
  IV U16902 ( .A(n17093), .Z(n17092) );
  XOR U16903 ( .A(n17094), .B(n17095), .Z(n17087) );
  ANDN U16904 ( .A(n17096), .B(n17039), .Z(n17095) );
  XNOR U16905 ( .A(n17094), .B(n17097), .Z(n17039) );
  XNOR U16906 ( .A(n17094), .B(n17037), .Z(n17096) );
  XOR U16907 ( .A(n17098), .B(n17099), .Z(n17037) );
  IV U16908 ( .A(n17100), .Z(n17099) );
  XOR U16909 ( .A(n17101), .B(n17102), .Z(n17094) );
  ANDN U16910 ( .A(n17103), .B(n17045), .Z(n17102) );
  XNOR U16911 ( .A(n17101), .B(n17104), .Z(n17045) );
  XNOR U16912 ( .A(n17101), .B(n17043), .Z(n17103) );
  XOR U16913 ( .A(n17105), .B(n17106), .Z(n17043) );
  IV U16914 ( .A(n17107), .Z(n17106) );
  XOR U16915 ( .A(n17108), .B(n17109), .Z(n17101) );
  NANDN U16916 ( .B(n17049), .A(n17110), .Z(n17108) );
  XOR U16917 ( .A(n17109), .B(n17047), .Z(n17110) );
  XOR U16918 ( .A(n17111), .B(n17112), .Z(n17047) );
  IV U16919 ( .A(n17113), .Z(n17112) );
  XNOR U16920 ( .A(n17114), .B(n17109), .Z(n17049) );
  OR U16921 ( .A(n11273), .B(n11274), .Z(n17109) );
  XOR U16922 ( .A(n17115), .B(n17116), .Z(n11273) );
  IV U16923 ( .A(n17117), .Z(n17116) );
  NAND U16924 ( .A(n16747), .B(n14945), .Z(n17114) );
  XOR U16925 ( .A(n16634), .B(n17118), .Z(n16627) );
  IV U16926 ( .A(n16633), .Z(n17118) );
  XNOR U16927 ( .A(n16630), .B(n17119), .Z(n16633) );
  XOR U16928 ( .A(n17120), .B(n17121), .Z(n16630) );
  ANDN U16929 ( .A(n17122), .B(n17058), .Z(n17121) );
  XNOR U16930 ( .A(n17120), .B(n17123), .Z(n17058) );
  XNOR U16931 ( .A(n17120), .B(n17056), .Z(n17122) );
  XOR U16932 ( .A(n17124), .B(n17125), .Z(n17056) );
  IV U16933 ( .A(n17126), .Z(n17125) );
  XOR U16934 ( .A(n17127), .B(n17128), .Z(n17120) );
  ANDN U16935 ( .A(n17129), .B(n17065), .Z(n17128) );
  XNOR U16936 ( .A(n17127), .B(n17130), .Z(n17065) );
  XNOR U16937 ( .A(n17127), .B(n17063), .Z(n17129) );
  XOR U16938 ( .A(n17131), .B(n17132), .Z(n17063) );
  IV U16939 ( .A(n17133), .Z(n17132) );
  XOR U16940 ( .A(n17134), .B(n17135), .Z(n17127) );
  ANDN U16941 ( .A(n17136), .B(n17072), .Z(n17135) );
  XNOR U16942 ( .A(n17134), .B(n17137), .Z(n17072) );
  XNOR U16943 ( .A(n17134), .B(n17070), .Z(n17136) );
  XOR U16944 ( .A(n17138), .B(n17139), .Z(n17070) );
  IV U16945 ( .A(n17140), .Z(n17139) );
  XOR U16946 ( .A(n17141), .B(n17142), .Z(n17134) );
  ANDN U16947 ( .A(n17143), .B(n17079), .Z(n17142) );
  XNOR U16948 ( .A(n17141), .B(n17144), .Z(n17079) );
  XNOR U16949 ( .A(n17141), .B(n17077), .Z(n17143) );
  XOR U16950 ( .A(n17145), .B(n17146), .Z(n17077) );
  IV U16951 ( .A(n17147), .Z(n17146) );
  XOR U16952 ( .A(n17148), .B(n17149), .Z(n17141) );
  ANDN U16953 ( .A(n17150), .B(n17086), .Z(n17149) );
  XNOR U16954 ( .A(n17148), .B(n17151), .Z(n17086) );
  XNOR U16955 ( .A(n17148), .B(n17084), .Z(n17150) );
  XOR U16956 ( .A(n17152), .B(n17153), .Z(n17084) );
  IV U16957 ( .A(n17154), .Z(n17153) );
  XOR U16958 ( .A(n17155), .B(n17156), .Z(n17148) );
  ANDN U16959 ( .A(n17157), .B(n17093), .Z(n17156) );
  XNOR U16960 ( .A(n17155), .B(n17158), .Z(n17093) );
  XNOR U16961 ( .A(n17155), .B(n17091), .Z(n17157) );
  XOR U16962 ( .A(n17159), .B(n17160), .Z(n17091) );
  IV U16963 ( .A(n17161), .Z(n17160) );
  XOR U16964 ( .A(n17162), .B(n17163), .Z(n17155) );
  ANDN U16965 ( .A(n17164), .B(n17100), .Z(n17163) );
  XNOR U16966 ( .A(n17162), .B(n17165), .Z(n17100) );
  XNOR U16967 ( .A(n17162), .B(n17098), .Z(n17164) );
  XOR U16968 ( .A(n17166), .B(n17167), .Z(n17098) );
  IV U16969 ( .A(n17168), .Z(n17167) );
  XOR U16970 ( .A(n17169), .B(n17170), .Z(n17162) );
  ANDN U16971 ( .A(n17171), .B(n17107), .Z(n17170) );
  XNOR U16972 ( .A(n17169), .B(n17172), .Z(n17107) );
  XNOR U16973 ( .A(n17169), .B(n17105), .Z(n17171) );
  XOR U16974 ( .A(n17173), .B(n17174), .Z(n17105) );
  IV U16975 ( .A(n17175), .Z(n17174) );
  XOR U16976 ( .A(n17176), .B(n17177), .Z(n17169) );
  ANDN U16977 ( .A(n17178), .B(n17113), .Z(n17177) );
  XNOR U16978 ( .A(n17176), .B(n17179), .Z(n17113) );
  XNOR U16979 ( .A(n17176), .B(n17111), .Z(n17178) );
  XOR U16980 ( .A(n17180), .B(n17181), .Z(n17111) );
  IV U16981 ( .A(n17182), .Z(n17181) );
  XOR U16982 ( .A(n17183), .B(n17184), .Z(n17176) );
  NANDN U16983 ( .B(n17117), .A(n17185), .Z(n17183) );
  XOR U16984 ( .A(n17184), .B(n17115), .Z(n17185) );
  XOR U16985 ( .A(n17186), .B(n17187), .Z(n17115) );
  IV U16986 ( .A(n17188), .Z(n17187) );
  XNOR U16987 ( .A(n17189), .B(n17184), .Z(n17117) );
  OR U16988 ( .A(n11413), .B(n11414), .Z(n17184) );
  XOR U16989 ( .A(n17190), .B(n17191), .Z(n11413) );
  IV U16990 ( .A(n17192), .Z(n17191) );
  NAND U16991 ( .A(n16747), .B(n15236), .Z(n17189) );
  XOR U16992 ( .A(n16641), .B(n17193), .Z(n16634) );
  IV U16993 ( .A(n16640), .Z(n17193) );
  XNOR U16994 ( .A(n16637), .B(n17194), .Z(n16640) );
  XOR U16995 ( .A(n17195), .B(n17196), .Z(n16637) );
  ANDN U16996 ( .A(n17197), .B(n17126), .Z(n17196) );
  XNOR U16997 ( .A(n17195), .B(n17198), .Z(n17126) );
  XNOR U16998 ( .A(n17195), .B(n17124), .Z(n17197) );
  XOR U16999 ( .A(n17199), .B(n17200), .Z(n17124) );
  IV U17000 ( .A(n17201), .Z(n17200) );
  XOR U17001 ( .A(n17202), .B(n17203), .Z(n17195) );
  ANDN U17002 ( .A(n17204), .B(n17133), .Z(n17203) );
  XNOR U17003 ( .A(n17202), .B(n17205), .Z(n17133) );
  XNOR U17004 ( .A(n17202), .B(n17131), .Z(n17204) );
  XOR U17005 ( .A(n17206), .B(n17207), .Z(n17131) );
  IV U17006 ( .A(n17208), .Z(n17207) );
  XOR U17007 ( .A(n17209), .B(n17210), .Z(n17202) );
  ANDN U17008 ( .A(n17211), .B(n17140), .Z(n17210) );
  XNOR U17009 ( .A(n17209), .B(n17212), .Z(n17140) );
  XNOR U17010 ( .A(n17209), .B(n17138), .Z(n17211) );
  XOR U17011 ( .A(n17213), .B(n17214), .Z(n17138) );
  IV U17012 ( .A(n17215), .Z(n17214) );
  XOR U17013 ( .A(n17216), .B(n17217), .Z(n17209) );
  ANDN U17014 ( .A(n17218), .B(n17147), .Z(n17217) );
  XNOR U17015 ( .A(n17216), .B(n17219), .Z(n17147) );
  XNOR U17016 ( .A(n17216), .B(n17145), .Z(n17218) );
  XOR U17017 ( .A(n17220), .B(n17221), .Z(n17145) );
  IV U17018 ( .A(n17222), .Z(n17221) );
  XOR U17019 ( .A(n17223), .B(n17224), .Z(n17216) );
  ANDN U17020 ( .A(n17225), .B(n17154), .Z(n17224) );
  XNOR U17021 ( .A(n17223), .B(n17226), .Z(n17154) );
  XNOR U17022 ( .A(n17223), .B(n17152), .Z(n17225) );
  XOR U17023 ( .A(n17227), .B(n17228), .Z(n17152) );
  IV U17024 ( .A(n17229), .Z(n17228) );
  XOR U17025 ( .A(n17230), .B(n17231), .Z(n17223) );
  ANDN U17026 ( .A(n17232), .B(n17161), .Z(n17231) );
  XNOR U17027 ( .A(n17230), .B(n17233), .Z(n17161) );
  XNOR U17028 ( .A(n17230), .B(n17159), .Z(n17232) );
  XOR U17029 ( .A(n17234), .B(n17235), .Z(n17159) );
  IV U17030 ( .A(n17236), .Z(n17235) );
  XOR U17031 ( .A(n17237), .B(n17238), .Z(n17230) );
  ANDN U17032 ( .A(n17239), .B(n17168), .Z(n17238) );
  XNOR U17033 ( .A(n17237), .B(n17240), .Z(n17168) );
  XNOR U17034 ( .A(n17237), .B(n17166), .Z(n17239) );
  XOR U17035 ( .A(n17241), .B(n17242), .Z(n17166) );
  IV U17036 ( .A(n17243), .Z(n17242) );
  XOR U17037 ( .A(n17244), .B(n17245), .Z(n17237) );
  ANDN U17038 ( .A(n17246), .B(n17175), .Z(n17245) );
  XNOR U17039 ( .A(n17244), .B(n17247), .Z(n17175) );
  XNOR U17040 ( .A(n17244), .B(n17173), .Z(n17246) );
  XOR U17041 ( .A(n17248), .B(n17249), .Z(n17173) );
  IV U17042 ( .A(n17250), .Z(n17249) );
  XOR U17043 ( .A(n17251), .B(n17252), .Z(n17244) );
  ANDN U17044 ( .A(n17253), .B(n17182), .Z(n17252) );
  XNOR U17045 ( .A(n17251), .B(n17254), .Z(n17182) );
  XNOR U17046 ( .A(n17251), .B(n17180), .Z(n17253) );
  XOR U17047 ( .A(n17255), .B(n17256), .Z(n17180) );
  IV U17048 ( .A(n17257), .Z(n17256) );
  XOR U17049 ( .A(n17258), .B(n17259), .Z(n17251) );
  ANDN U17050 ( .A(n17260), .B(n17188), .Z(n17259) );
  XNOR U17051 ( .A(n17258), .B(n17261), .Z(n17188) );
  XNOR U17052 ( .A(n17258), .B(n17186), .Z(n17260) );
  XOR U17053 ( .A(n17262), .B(n17263), .Z(n17186) );
  IV U17054 ( .A(n17264), .Z(n17263) );
  XOR U17055 ( .A(n17265), .B(n17266), .Z(n17258) );
  NANDN U17056 ( .B(n17192), .A(n17267), .Z(n17265) );
  XOR U17057 ( .A(n17266), .B(n17190), .Z(n17267) );
  XOR U17058 ( .A(n17268), .B(n17269), .Z(n17190) );
  IV U17059 ( .A(n17270), .Z(n17269) );
  XNOR U17060 ( .A(n17271), .B(n17266), .Z(n17192) );
  OR U17061 ( .A(n11546), .B(n11547), .Z(n17266) );
  XOR U17062 ( .A(n17272), .B(n17273), .Z(n11546) );
  IV U17063 ( .A(n17274), .Z(n17273) );
  NAND U17064 ( .A(n16747), .B(n15553), .Z(n17271) );
  XOR U17065 ( .A(n16648), .B(n17275), .Z(n16641) );
  IV U17066 ( .A(n16647), .Z(n17275) );
  XNOR U17067 ( .A(n16644), .B(n17276), .Z(n16647) );
  XOR U17068 ( .A(n17277), .B(n17278), .Z(n16644) );
  ANDN U17069 ( .A(n17279), .B(n17201), .Z(n17278) );
  XNOR U17070 ( .A(n17277), .B(n17280), .Z(n17201) );
  XNOR U17071 ( .A(n17277), .B(n17199), .Z(n17279) );
  XOR U17072 ( .A(n17281), .B(n17282), .Z(n17199) );
  IV U17073 ( .A(n17283), .Z(n17282) );
  XOR U17074 ( .A(n17284), .B(n17285), .Z(n17277) );
  ANDN U17075 ( .A(n17286), .B(n17208), .Z(n17285) );
  XNOR U17076 ( .A(n17284), .B(n17287), .Z(n17208) );
  XNOR U17077 ( .A(n17284), .B(n17206), .Z(n17286) );
  XOR U17078 ( .A(n17288), .B(n17289), .Z(n17206) );
  IV U17079 ( .A(n17290), .Z(n17289) );
  XOR U17080 ( .A(n17291), .B(n17292), .Z(n17284) );
  ANDN U17081 ( .A(n17293), .B(n17215), .Z(n17292) );
  XNOR U17082 ( .A(n17291), .B(n17294), .Z(n17215) );
  XNOR U17083 ( .A(n17291), .B(n17213), .Z(n17293) );
  XOR U17084 ( .A(n17295), .B(n17296), .Z(n17213) );
  IV U17085 ( .A(n17297), .Z(n17296) );
  XOR U17086 ( .A(n17298), .B(n17299), .Z(n17291) );
  ANDN U17087 ( .A(n17300), .B(n17222), .Z(n17299) );
  XNOR U17088 ( .A(n17298), .B(n17301), .Z(n17222) );
  XNOR U17089 ( .A(n17298), .B(n17220), .Z(n17300) );
  XOR U17090 ( .A(n17302), .B(n17303), .Z(n17220) );
  IV U17091 ( .A(n17304), .Z(n17303) );
  XOR U17092 ( .A(n17305), .B(n17306), .Z(n17298) );
  ANDN U17093 ( .A(n17307), .B(n17229), .Z(n17306) );
  XNOR U17094 ( .A(n17305), .B(n17308), .Z(n17229) );
  XNOR U17095 ( .A(n17305), .B(n17227), .Z(n17307) );
  XOR U17096 ( .A(n17309), .B(n17310), .Z(n17227) );
  IV U17097 ( .A(n17311), .Z(n17310) );
  XOR U17098 ( .A(n17312), .B(n17313), .Z(n17305) );
  ANDN U17099 ( .A(n17314), .B(n17236), .Z(n17313) );
  XNOR U17100 ( .A(n17312), .B(n17315), .Z(n17236) );
  XNOR U17101 ( .A(n17312), .B(n17234), .Z(n17314) );
  XOR U17102 ( .A(n17316), .B(n17317), .Z(n17234) );
  IV U17103 ( .A(n17318), .Z(n17317) );
  XOR U17104 ( .A(n17319), .B(n17320), .Z(n17312) );
  ANDN U17105 ( .A(n17321), .B(n17243), .Z(n17320) );
  XNOR U17106 ( .A(n17319), .B(n17322), .Z(n17243) );
  XNOR U17107 ( .A(n17319), .B(n17241), .Z(n17321) );
  XOR U17108 ( .A(n17323), .B(n17324), .Z(n17241) );
  IV U17109 ( .A(n17325), .Z(n17324) );
  XOR U17110 ( .A(n17326), .B(n17327), .Z(n17319) );
  ANDN U17111 ( .A(n17328), .B(n17250), .Z(n17327) );
  XNOR U17112 ( .A(n17326), .B(n17329), .Z(n17250) );
  XNOR U17113 ( .A(n17326), .B(n17248), .Z(n17328) );
  XOR U17114 ( .A(n17330), .B(n17331), .Z(n17248) );
  IV U17115 ( .A(n17332), .Z(n17331) );
  XOR U17116 ( .A(n17333), .B(n17334), .Z(n17326) );
  ANDN U17117 ( .A(n17335), .B(n17257), .Z(n17334) );
  XNOR U17118 ( .A(n17333), .B(n17336), .Z(n17257) );
  XNOR U17119 ( .A(n17333), .B(n17255), .Z(n17335) );
  XOR U17120 ( .A(n17337), .B(n17338), .Z(n17255) );
  IV U17121 ( .A(n17339), .Z(n17338) );
  XOR U17122 ( .A(n17340), .B(n17341), .Z(n17333) );
  ANDN U17123 ( .A(n17342), .B(n17264), .Z(n17341) );
  XNOR U17124 ( .A(n17340), .B(n17343), .Z(n17264) );
  XNOR U17125 ( .A(n17340), .B(n17262), .Z(n17342) );
  XOR U17126 ( .A(n17344), .B(n17345), .Z(n17262) );
  IV U17127 ( .A(n17346), .Z(n17345) );
  XOR U17128 ( .A(n17347), .B(n17348), .Z(n17340) );
  ANDN U17129 ( .A(n17349), .B(n17270), .Z(n17348) );
  XNOR U17130 ( .A(n17347), .B(n17350), .Z(n17270) );
  XNOR U17131 ( .A(n17347), .B(n17268), .Z(n17349) );
  XOR U17132 ( .A(n17351), .B(n17352), .Z(n17268) );
  IV U17133 ( .A(n17353), .Z(n17352) );
  XOR U17134 ( .A(n17354), .B(n17355), .Z(n17347) );
  NANDN U17135 ( .B(n17274), .A(n17356), .Z(n17354) );
  XOR U17136 ( .A(n17355), .B(n17272), .Z(n17356) );
  XOR U17137 ( .A(n17357), .B(n17358), .Z(n17272) );
  IV U17138 ( .A(n17359), .Z(n17358) );
  XNOR U17139 ( .A(n17360), .B(n17355), .Z(n17274) );
  OR U17140 ( .A(n11673), .B(n11674), .Z(n17355) );
  XOR U17141 ( .A(n17361), .B(n17362), .Z(n11673) );
  IV U17142 ( .A(n17363), .Z(n17362) );
  NAND U17143 ( .A(n16747), .B(n15896), .Z(n17360) );
  XOR U17144 ( .A(n16655), .B(n17364), .Z(n16648) );
  IV U17145 ( .A(n16654), .Z(n17364) );
  XNOR U17146 ( .A(n16651), .B(n17365), .Z(n16654) );
  XOR U17147 ( .A(n17366), .B(n17367), .Z(n16651) );
  ANDN U17148 ( .A(n17368), .B(n17283), .Z(n17367) );
  XNOR U17149 ( .A(n17366), .B(n17369), .Z(n17283) );
  XNOR U17150 ( .A(n17366), .B(n17281), .Z(n17368) );
  XOR U17151 ( .A(n17370), .B(n17371), .Z(n17281) );
  IV U17152 ( .A(n17372), .Z(n17371) );
  XOR U17153 ( .A(n17373), .B(n17374), .Z(n17366) );
  ANDN U17154 ( .A(n17375), .B(n17290), .Z(n17374) );
  XNOR U17155 ( .A(n17373), .B(n17376), .Z(n17290) );
  XNOR U17156 ( .A(n17373), .B(n17288), .Z(n17375) );
  XOR U17157 ( .A(n17377), .B(n17378), .Z(n17288) );
  IV U17158 ( .A(n17379), .Z(n17378) );
  XOR U17159 ( .A(n17380), .B(n17381), .Z(n17373) );
  ANDN U17160 ( .A(n17382), .B(n17297), .Z(n17381) );
  XNOR U17161 ( .A(n17380), .B(n17383), .Z(n17297) );
  XNOR U17162 ( .A(n17380), .B(n17295), .Z(n17382) );
  XOR U17163 ( .A(n17384), .B(n17385), .Z(n17295) );
  IV U17164 ( .A(n17386), .Z(n17385) );
  XOR U17165 ( .A(n17387), .B(n17388), .Z(n17380) );
  ANDN U17166 ( .A(n17389), .B(n17304), .Z(n17388) );
  XNOR U17167 ( .A(n17387), .B(n17390), .Z(n17304) );
  XNOR U17168 ( .A(n17387), .B(n17302), .Z(n17389) );
  XOR U17169 ( .A(n17391), .B(n17392), .Z(n17302) );
  IV U17170 ( .A(n17393), .Z(n17392) );
  XOR U17171 ( .A(n17394), .B(n17395), .Z(n17387) );
  ANDN U17172 ( .A(n17396), .B(n17311), .Z(n17395) );
  XNOR U17173 ( .A(n17394), .B(n17397), .Z(n17311) );
  XNOR U17174 ( .A(n17394), .B(n17309), .Z(n17396) );
  XOR U17175 ( .A(n17398), .B(n17399), .Z(n17309) );
  IV U17176 ( .A(n17400), .Z(n17399) );
  XOR U17177 ( .A(n17401), .B(n17402), .Z(n17394) );
  ANDN U17178 ( .A(n17403), .B(n17318), .Z(n17402) );
  XNOR U17179 ( .A(n17401), .B(n17404), .Z(n17318) );
  XNOR U17180 ( .A(n17401), .B(n17316), .Z(n17403) );
  XOR U17181 ( .A(n17405), .B(n17406), .Z(n17316) );
  IV U17182 ( .A(n17407), .Z(n17406) );
  XOR U17183 ( .A(n17408), .B(n17409), .Z(n17401) );
  ANDN U17184 ( .A(n17410), .B(n17325), .Z(n17409) );
  XNOR U17185 ( .A(n17408), .B(n17411), .Z(n17325) );
  XNOR U17186 ( .A(n17408), .B(n17323), .Z(n17410) );
  XOR U17187 ( .A(n17412), .B(n17413), .Z(n17323) );
  IV U17188 ( .A(n17414), .Z(n17413) );
  XOR U17189 ( .A(n17415), .B(n17416), .Z(n17408) );
  ANDN U17190 ( .A(n17417), .B(n17332), .Z(n17416) );
  XNOR U17191 ( .A(n17415), .B(n17418), .Z(n17332) );
  XNOR U17192 ( .A(n17415), .B(n17330), .Z(n17417) );
  XOR U17193 ( .A(n17419), .B(n17420), .Z(n17330) );
  IV U17194 ( .A(n17421), .Z(n17420) );
  XOR U17195 ( .A(n17422), .B(n17423), .Z(n17415) );
  ANDN U17196 ( .A(n17424), .B(n17339), .Z(n17423) );
  XNOR U17197 ( .A(n17422), .B(n17425), .Z(n17339) );
  XNOR U17198 ( .A(n17422), .B(n17337), .Z(n17424) );
  XOR U17199 ( .A(n17426), .B(n17427), .Z(n17337) );
  IV U17200 ( .A(n17428), .Z(n17427) );
  XOR U17201 ( .A(n17429), .B(n17430), .Z(n17422) );
  ANDN U17202 ( .A(n17431), .B(n17346), .Z(n17430) );
  XNOR U17203 ( .A(n17429), .B(n17432), .Z(n17346) );
  XNOR U17204 ( .A(n17429), .B(n17344), .Z(n17431) );
  XOR U17205 ( .A(n17433), .B(n17434), .Z(n17344) );
  IV U17206 ( .A(n17435), .Z(n17434) );
  XOR U17207 ( .A(n17436), .B(n17437), .Z(n17429) );
  ANDN U17208 ( .A(n17438), .B(n17353), .Z(n17437) );
  XNOR U17209 ( .A(n17436), .B(n17439), .Z(n17353) );
  XNOR U17210 ( .A(n17436), .B(n17351), .Z(n17438) );
  XOR U17211 ( .A(n17440), .B(n17441), .Z(n17351) );
  IV U17212 ( .A(n17442), .Z(n17441) );
  XOR U17213 ( .A(n17443), .B(n17444), .Z(n17436) );
  ANDN U17214 ( .A(n17445), .B(n17359), .Z(n17444) );
  XNOR U17215 ( .A(n17443), .B(n17446), .Z(n17359) );
  XNOR U17216 ( .A(n17443), .B(n17357), .Z(n17445) );
  XOR U17217 ( .A(n17447), .B(n17448), .Z(n17357) );
  IV U17218 ( .A(n17449), .Z(n17448) );
  XOR U17219 ( .A(n17450), .B(n17451), .Z(n17443) );
  NANDN U17220 ( .B(n17363), .A(n17452), .Z(n17450) );
  XOR U17221 ( .A(n17451), .B(n17361), .Z(n17452) );
  XOR U17222 ( .A(n17453), .B(n17454), .Z(n17361) );
  IV U17223 ( .A(n17455), .Z(n17454) );
  XNOR U17224 ( .A(n17456), .B(n17451), .Z(n17363) );
  OR U17225 ( .A(n11686), .B(n11687), .Z(n17451) );
  XOR U17226 ( .A(n17457), .B(n17458), .Z(n11686) );
  IV U17227 ( .A(n17459), .Z(n17458) );
  NAND U17228 ( .A(n16747), .B(n16265), .Z(n17456) );
  XOR U17229 ( .A(n16662), .B(n17460), .Z(n16655) );
  IV U17230 ( .A(n16661), .Z(n17460) );
  XNOR U17231 ( .A(n16658), .B(n17461), .Z(n16661) );
  XOR U17232 ( .A(n17462), .B(n17463), .Z(n16658) );
  ANDN U17233 ( .A(n17464), .B(n17372), .Z(n17463) );
  XNOR U17234 ( .A(n17462), .B(n17465), .Z(n17372) );
  XNOR U17235 ( .A(n17462), .B(n17370), .Z(n17464) );
  XOR U17236 ( .A(n17466), .B(n17467), .Z(n17370) );
  IV U17237 ( .A(n17468), .Z(n17467) );
  XOR U17238 ( .A(n17469), .B(n17470), .Z(n17462) );
  ANDN U17239 ( .A(n17471), .B(n17379), .Z(n17470) );
  XNOR U17240 ( .A(n17469), .B(n17472), .Z(n17379) );
  XNOR U17241 ( .A(n17469), .B(n17377), .Z(n17471) );
  XOR U17242 ( .A(n17473), .B(n17474), .Z(n17377) );
  IV U17243 ( .A(n17475), .Z(n17474) );
  XOR U17244 ( .A(n17476), .B(n17477), .Z(n17469) );
  ANDN U17245 ( .A(n17478), .B(n17386), .Z(n17477) );
  XNOR U17246 ( .A(n17476), .B(n17479), .Z(n17386) );
  XNOR U17247 ( .A(n17476), .B(n17384), .Z(n17478) );
  XOR U17248 ( .A(n17480), .B(n17481), .Z(n17384) );
  IV U17249 ( .A(n17482), .Z(n17481) );
  XOR U17250 ( .A(n17483), .B(n17484), .Z(n17476) );
  ANDN U17251 ( .A(n17485), .B(n17393), .Z(n17484) );
  XNOR U17252 ( .A(n17483), .B(n17486), .Z(n17393) );
  XNOR U17253 ( .A(n17483), .B(n17391), .Z(n17485) );
  XOR U17254 ( .A(n17487), .B(n17488), .Z(n17391) );
  IV U17255 ( .A(n17489), .Z(n17488) );
  XOR U17256 ( .A(n17490), .B(n17491), .Z(n17483) );
  ANDN U17257 ( .A(n17492), .B(n17400), .Z(n17491) );
  XNOR U17258 ( .A(n17490), .B(n17493), .Z(n17400) );
  XNOR U17259 ( .A(n17490), .B(n17398), .Z(n17492) );
  XOR U17260 ( .A(n17494), .B(n17495), .Z(n17398) );
  IV U17261 ( .A(n17496), .Z(n17495) );
  XOR U17262 ( .A(n17497), .B(n17498), .Z(n17490) );
  ANDN U17263 ( .A(n17499), .B(n17407), .Z(n17498) );
  XNOR U17264 ( .A(n17497), .B(n17500), .Z(n17407) );
  XNOR U17265 ( .A(n17497), .B(n17405), .Z(n17499) );
  XOR U17266 ( .A(n17501), .B(n17502), .Z(n17405) );
  IV U17267 ( .A(n17503), .Z(n17502) );
  XOR U17268 ( .A(n17504), .B(n17505), .Z(n17497) );
  ANDN U17269 ( .A(n17506), .B(n17414), .Z(n17505) );
  XNOR U17270 ( .A(n17504), .B(n17507), .Z(n17414) );
  XNOR U17271 ( .A(n17504), .B(n17412), .Z(n17506) );
  XOR U17272 ( .A(n17508), .B(n17509), .Z(n17412) );
  IV U17273 ( .A(n17510), .Z(n17509) );
  XOR U17274 ( .A(n17511), .B(n17512), .Z(n17504) );
  ANDN U17275 ( .A(n17513), .B(n17421), .Z(n17512) );
  XNOR U17276 ( .A(n17511), .B(n17514), .Z(n17421) );
  XNOR U17277 ( .A(n17511), .B(n17419), .Z(n17513) );
  XOR U17278 ( .A(n17515), .B(n17516), .Z(n17419) );
  IV U17279 ( .A(n17517), .Z(n17516) );
  XOR U17280 ( .A(n17518), .B(n17519), .Z(n17511) );
  ANDN U17281 ( .A(n17520), .B(n17428), .Z(n17519) );
  XNOR U17282 ( .A(n17518), .B(n17521), .Z(n17428) );
  XNOR U17283 ( .A(n17518), .B(n17426), .Z(n17520) );
  XOR U17284 ( .A(n17522), .B(n17523), .Z(n17426) );
  IV U17285 ( .A(n17524), .Z(n17523) );
  XOR U17286 ( .A(n17525), .B(n17526), .Z(n17518) );
  ANDN U17287 ( .A(n17527), .B(n17435), .Z(n17526) );
  XNOR U17288 ( .A(n17525), .B(n17528), .Z(n17435) );
  XNOR U17289 ( .A(n17525), .B(n17433), .Z(n17527) );
  XOR U17290 ( .A(n17529), .B(n17530), .Z(n17433) );
  IV U17291 ( .A(n17531), .Z(n17530) );
  XOR U17292 ( .A(n17532), .B(n17533), .Z(n17525) );
  ANDN U17293 ( .A(n17534), .B(n17442), .Z(n17533) );
  XNOR U17294 ( .A(n17532), .B(n17535), .Z(n17442) );
  XNOR U17295 ( .A(n17532), .B(n17440), .Z(n17534) );
  XOR U17296 ( .A(n17536), .B(n17537), .Z(n17440) );
  IV U17297 ( .A(n17538), .Z(n17537) );
  XOR U17298 ( .A(n17539), .B(n17540), .Z(n17532) );
  ANDN U17299 ( .A(n17541), .B(n17449), .Z(n17540) );
  XNOR U17300 ( .A(n17539), .B(n17542), .Z(n17449) );
  XNOR U17301 ( .A(n17539), .B(n17447), .Z(n17541) );
  XOR U17302 ( .A(n17543), .B(n17544), .Z(n17447) );
  IV U17303 ( .A(n17545), .Z(n17544) );
  XOR U17304 ( .A(n17546), .B(n17547), .Z(n17539) );
  ANDN U17305 ( .A(n17548), .B(n17455), .Z(n17547) );
  XNOR U17306 ( .A(n17546), .B(n17549), .Z(n17455) );
  XNOR U17307 ( .A(n17546), .B(n17453), .Z(n17548) );
  XOR U17308 ( .A(n17550), .B(n17551), .Z(n17453) );
  IV U17309 ( .A(n17552), .Z(n17551) );
  XOR U17310 ( .A(n17553), .B(n17554), .Z(n17546) );
  NANDN U17311 ( .B(n17459), .A(n17555), .Z(n17553) );
  XOR U17312 ( .A(n17554), .B(n17457), .Z(n17555) );
  XOR U17313 ( .A(n17556), .B(n17557), .Z(n17457) );
  IV U17314 ( .A(n17558), .Z(n17557) );
  XNOR U17315 ( .A(n17559), .B(n17554), .Z(n17459) );
  OR U17316 ( .A(n11819), .B(n11820), .Z(n17554) );
  XOR U17317 ( .A(n17560), .B(n17561), .Z(n11819) );
  IV U17318 ( .A(n17562), .Z(n17561) );
  NAND U17319 ( .A(n16747), .B(n16657), .Z(n17559) );
  XOR U17320 ( .A(n16668), .B(n17563), .Z(n16662) );
  IV U17321 ( .A(n16667), .Z(n17563) );
  XNOR U17322 ( .A(n16664), .B(n17461), .Z(n16667) );
  AND U17323 ( .A(n17567), .B(n16657), .Z(n17461) );
  XOR U17324 ( .A(n17564), .B(n17565), .Z(n16664) );
  ANDN U17325 ( .A(n17566), .B(n17468), .Z(n17565) );
  XNOR U17326 ( .A(n17564), .B(n17567), .Z(n17468) );
  XNOR U17327 ( .A(n17564), .B(n17466), .Z(n17566) );
  XOR U17328 ( .A(n17568), .B(n17569), .Z(n17466) );
  IV U17329 ( .A(n17570), .Z(n17569) );
  XOR U17330 ( .A(n17571), .B(n17572), .Z(n17564) );
  ANDN U17331 ( .A(n17573), .B(n17475), .Z(n17572) );
  XNOR U17332 ( .A(n17571), .B(n17574), .Z(n17475) );
  XNOR U17333 ( .A(n17571), .B(n17473), .Z(n17573) );
  XOR U17334 ( .A(n17575), .B(n17576), .Z(n17473) );
  IV U17335 ( .A(n17577), .Z(n17576) );
  XOR U17336 ( .A(n17578), .B(n17579), .Z(n17571) );
  ANDN U17337 ( .A(n17580), .B(n17482), .Z(n17579) );
  XNOR U17338 ( .A(n17578), .B(n17581), .Z(n17482) );
  XNOR U17339 ( .A(n17578), .B(n17480), .Z(n17580) );
  XOR U17340 ( .A(n17582), .B(n17583), .Z(n17480) );
  IV U17341 ( .A(n17584), .Z(n17583) );
  XOR U17342 ( .A(n17585), .B(n17586), .Z(n17578) );
  ANDN U17343 ( .A(n17587), .B(n17489), .Z(n17586) );
  XNOR U17344 ( .A(n17585), .B(n17588), .Z(n17489) );
  XNOR U17345 ( .A(n17585), .B(n17487), .Z(n17587) );
  XOR U17346 ( .A(n17589), .B(n17590), .Z(n17487) );
  IV U17347 ( .A(n17591), .Z(n17590) );
  XOR U17348 ( .A(n17592), .B(n17593), .Z(n17585) );
  ANDN U17349 ( .A(n17594), .B(n17496), .Z(n17593) );
  XNOR U17350 ( .A(n17592), .B(n17595), .Z(n17496) );
  XNOR U17351 ( .A(n17592), .B(n17494), .Z(n17594) );
  XOR U17352 ( .A(n17596), .B(n17597), .Z(n17494) );
  IV U17353 ( .A(n17598), .Z(n17597) );
  XOR U17354 ( .A(n17599), .B(n17600), .Z(n17592) );
  ANDN U17355 ( .A(n17601), .B(n17503), .Z(n17600) );
  XNOR U17356 ( .A(n17599), .B(n17602), .Z(n17503) );
  XNOR U17357 ( .A(n17599), .B(n17501), .Z(n17601) );
  XOR U17358 ( .A(n17603), .B(n17604), .Z(n17501) );
  IV U17359 ( .A(n17605), .Z(n17604) );
  XOR U17360 ( .A(n17606), .B(n17607), .Z(n17599) );
  ANDN U17361 ( .A(n17608), .B(n17510), .Z(n17607) );
  XNOR U17362 ( .A(n17606), .B(n17609), .Z(n17510) );
  XNOR U17363 ( .A(n17606), .B(n17508), .Z(n17608) );
  XOR U17364 ( .A(n17610), .B(n17611), .Z(n17508) );
  IV U17365 ( .A(n17612), .Z(n17611) );
  XOR U17366 ( .A(n17613), .B(n17614), .Z(n17606) );
  ANDN U17367 ( .A(n17615), .B(n17517), .Z(n17614) );
  XNOR U17368 ( .A(n17613), .B(n17616), .Z(n17517) );
  XNOR U17369 ( .A(n17613), .B(n17515), .Z(n17615) );
  XOR U17370 ( .A(n17617), .B(n17618), .Z(n17515) );
  IV U17371 ( .A(n17619), .Z(n17618) );
  XOR U17372 ( .A(n17620), .B(n17621), .Z(n17613) );
  ANDN U17373 ( .A(n17622), .B(n17524), .Z(n17621) );
  XNOR U17374 ( .A(n17620), .B(n17623), .Z(n17524) );
  XNOR U17375 ( .A(n17620), .B(n17522), .Z(n17622) );
  XOR U17376 ( .A(n17624), .B(n17625), .Z(n17522) );
  IV U17377 ( .A(n17626), .Z(n17625) );
  XOR U17378 ( .A(n17627), .B(n17628), .Z(n17620) );
  ANDN U17379 ( .A(n17629), .B(n17531), .Z(n17628) );
  XNOR U17380 ( .A(n17627), .B(n17630), .Z(n17531) );
  XNOR U17381 ( .A(n17627), .B(n17529), .Z(n17629) );
  XOR U17382 ( .A(n17631), .B(n17632), .Z(n17529) );
  IV U17383 ( .A(n17633), .Z(n17632) );
  XOR U17384 ( .A(n17634), .B(n17635), .Z(n17627) );
  ANDN U17385 ( .A(n17636), .B(n17538), .Z(n17635) );
  XNOR U17386 ( .A(n17634), .B(n17637), .Z(n17538) );
  XNOR U17387 ( .A(n17634), .B(n17536), .Z(n17636) );
  XOR U17388 ( .A(n17638), .B(n17639), .Z(n17536) );
  IV U17389 ( .A(n17640), .Z(n17639) );
  XOR U17390 ( .A(n17641), .B(n17642), .Z(n17634) );
  ANDN U17391 ( .A(n17643), .B(n17545), .Z(n17642) );
  XNOR U17392 ( .A(n17641), .B(n17644), .Z(n17545) );
  XNOR U17393 ( .A(n17641), .B(n17543), .Z(n17643) );
  XOR U17394 ( .A(n17645), .B(n17646), .Z(n17543) );
  IV U17395 ( .A(n17647), .Z(n17646) );
  XOR U17396 ( .A(n17648), .B(n17649), .Z(n17641) );
  ANDN U17397 ( .A(n17650), .B(n17552), .Z(n17649) );
  XNOR U17398 ( .A(n17648), .B(n17651), .Z(n17552) );
  XNOR U17399 ( .A(n17648), .B(n17550), .Z(n17650) );
  XOR U17400 ( .A(n17652), .B(n17653), .Z(n17550) );
  IV U17401 ( .A(n17654), .Z(n17653) );
  XOR U17402 ( .A(n17655), .B(n17656), .Z(n17648) );
  ANDN U17403 ( .A(n17657), .B(n17558), .Z(n17656) );
  XNOR U17404 ( .A(n17655), .B(n17658), .Z(n17558) );
  XNOR U17405 ( .A(n17655), .B(n17556), .Z(n17657) );
  XOR U17406 ( .A(n17659), .B(n17660), .Z(n17556) );
  IV U17407 ( .A(n17661), .Z(n17660) );
  XOR U17408 ( .A(n17662), .B(n17663), .Z(n17655) );
  NANDN U17409 ( .B(n17562), .A(n17664), .Z(n17662) );
  XOR U17410 ( .A(n17663), .B(n17560), .Z(n17664) );
  XOR U17411 ( .A(n17665), .B(n17666), .Z(n17560) );
  IV U17412 ( .A(n17667), .Z(n17666) );
  XNOR U17413 ( .A(n17668), .B(n17663), .Z(n17562) );
  OR U17414 ( .A(n11952), .B(n11953), .Z(n17663) );
  XOR U17415 ( .A(n17669), .B(n17670), .Z(n11952) );
  IV U17416 ( .A(n17671), .Z(n17670) );
  NAND U17417 ( .A(n16747), .B(n17567), .Z(n17668) );
  XOR U17418 ( .A(n16674), .B(n17672), .Z(n16668) );
  IV U17419 ( .A(n16673), .Z(n17672) );
  XNOR U17420 ( .A(n16670), .B(n17365), .Z(n16673) );
  AND U17421 ( .A(n17688), .B(n16265), .Z(n17365) );
  XOR U17422 ( .A(n17673), .B(n17674), .Z(n16670) );
  ANDN U17423 ( .A(n17675), .B(n17570), .Z(n17674) );
  XNOR U17424 ( .A(n17673), .B(n17465), .Z(n17570) );
  AND U17425 ( .A(n17688), .B(n16657), .Z(n17465) );
  XNOR U17426 ( .A(n17673), .B(n17568), .Z(n17675) );
  XOR U17427 ( .A(n17676), .B(n17677), .Z(n17568) );
  IV U17428 ( .A(n17678), .Z(n17677) );
  XOR U17429 ( .A(n17679), .B(n17680), .Z(n17673) );
  ANDN U17430 ( .A(n17681), .B(n17577), .Z(n17680) );
  XNOR U17431 ( .A(n17679), .B(n17574), .Z(n17577) );
  AND U17432 ( .A(n17688), .B(n17567), .Z(n17574) );
  XNOR U17433 ( .A(n17679), .B(n17575), .Z(n17681) );
  XOR U17434 ( .A(n17682), .B(n17683), .Z(n17575) );
  IV U17435 ( .A(n17684), .Z(n17683) );
  XOR U17436 ( .A(n17685), .B(n17686), .Z(n17679) );
  ANDN U17437 ( .A(n17687), .B(n17584), .Z(n17686) );
  XNOR U17438 ( .A(n17685), .B(n17688), .Z(n17584) );
  XNOR U17439 ( .A(n17685), .B(n17582), .Z(n17687) );
  XOR U17440 ( .A(n17689), .B(n17690), .Z(n17582) );
  IV U17441 ( .A(n17691), .Z(n17690) );
  XOR U17442 ( .A(n17692), .B(n17693), .Z(n17685) );
  ANDN U17443 ( .A(n17694), .B(n17591), .Z(n17693) );
  XNOR U17444 ( .A(n17692), .B(n17695), .Z(n17591) );
  XNOR U17445 ( .A(n17692), .B(n17589), .Z(n17694) );
  XOR U17446 ( .A(n17696), .B(n17697), .Z(n17589) );
  IV U17447 ( .A(n17698), .Z(n17697) );
  XOR U17448 ( .A(n17699), .B(n17700), .Z(n17692) );
  ANDN U17449 ( .A(n17701), .B(n17598), .Z(n17700) );
  XNOR U17450 ( .A(n17699), .B(n17702), .Z(n17598) );
  XNOR U17451 ( .A(n17699), .B(n17596), .Z(n17701) );
  XOR U17452 ( .A(n17703), .B(n17704), .Z(n17596) );
  IV U17453 ( .A(n17705), .Z(n17704) );
  XOR U17454 ( .A(n17706), .B(n17707), .Z(n17699) );
  ANDN U17455 ( .A(n17708), .B(n17605), .Z(n17707) );
  XNOR U17456 ( .A(n17706), .B(n17709), .Z(n17605) );
  XNOR U17457 ( .A(n17706), .B(n17603), .Z(n17708) );
  XOR U17458 ( .A(n17710), .B(n17711), .Z(n17603) );
  IV U17459 ( .A(n17712), .Z(n17711) );
  XOR U17460 ( .A(n17713), .B(n17714), .Z(n17706) );
  ANDN U17461 ( .A(n17715), .B(n17612), .Z(n17714) );
  XNOR U17462 ( .A(n17713), .B(n17716), .Z(n17612) );
  XNOR U17463 ( .A(n17713), .B(n17610), .Z(n17715) );
  XOR U17464 ( .A(n17717), .B(n17718), .Z(n17610) );
  IV U17465 ( .A(n17719), .Z(n17718) );
  XOR U17466 ( .A(n17720), .B(n17721), .Z(n17713) );
  ANDN U17467 ( .A(n17722), .B(n17619), .Z(n17721) );
  XNOR U17468 ( .A(n17720), .B(n17723), .Z(n17619) );
  XNOR U17469 ( .A(n17720), .B(n17617), .Z(n17722) );
  XOR U17470 ( .A(n17724), .B(n17725), .Z(n17617) );
  IV U17471 ( .A(n17726), .Z(n17725) );
  XOR U17472 ( .A(n17727), .B(n17728), .Z(n17720) );
  ANDN U17473 ( .A(n17729), .B(n17626), .Z(n17728) );
  XNOR U17474 ( .A(n17727), .B(n17730), .Z(n17626) );
  XNOR U17475 ( .A(n17727), .B(n17624), .Z(n17729) );
  XOR U17476 ( .A(n17731), .B(n17732), .Z(n17624) );
  IV U17477 ( .A(n17733), .Z(n17732) );
  XOR U17478 ( .A(n17734), .B(n17735), .Z(n17727) );
  ANDN U17479 ( .A(n17736), .B(n17633), .Z(n17735) );
  XNOR U17480 ( .A(n17734), .B(n17737), .Z(n17633) );
  XNOR U17481 ( .A(n17734), .B(n17631), .Z(n17736) );
  XOR U17482 ( .A(n17738), .B(n17739), .Z(n17631) );
  IV U17483 ( .A(n17740), .Z(n17739) );
  XOR U17484 ( .A(n17741), .B(n17742), .Z(n17734) );
  ANDN U17485 ( .A(n17743), .B(n17640), .Z(n17742) );
  XNOR U17486 ( .A(n17741), .B(n17744), .Z(n17640) );
  XNOR U17487 ( .A(n17741), .B(n17638), .Z(n17743) );
  XOR U17488 ( .A(n17745), .B(n17746), .Z(n17638) );
  IV U17489 ( .A(n17747), .Z(n17746) );
  XOR U17490 ( .A(n17748), .B(n17749), .Z(n17741) );
  ANDN U17491 ( .A(n17750), .B(n17647), .Z(n17749) );
  XNOR U17492 ( .A(n17748), .B(n17751), .Z(n17647) );
  XNOR U17493 ( .A(n17748), .B(n17645), .Z(n17750) );
  XOR U17494 ( .A(n17752), .B(n17753), .Z(n17645) );
  IV U17495 ( .A(n17754), .Z(n17753) );
  XOR U17496 ( .A(n17755), .B(n17756), .Z(n17748) );
  ANDN U17497 ( .A(n17757), .B(n17654), .Z(n17756) );
  XNOR U17498 ( .A(n17755), .B(n17758), .Z(n17654) );
  XNOR U17499 ( .A(n17755), .B(n17652), .Z(n17757) );
  XOR U17500 ( .A(n17759), .B(n17760), .Z(n17652) );
  IV U17501 ( .A(n17761), .Z(n17760) );
  XOR U17502 ( .A(n17762), .B(n17763), .Z(n17755) );
  ANDN U17503 ( .A(n17764), .B(n17661), .Z(n17763) );
  XNOR U17504 ( .A(n17762), .B(n17765), .Z(n17661) );
  XNOR U17505 ( .A(n17762), .B(n17659), .Z(n17764) );
  XOR U17506 ( .A(n17766), .B(n17767), .Z(n17659) );
  IV U17507 ( .A(n17768), .Z(n17767) );
  XOR U17508 ( .A(n17769), .B(n17770), .Z(n17762) );
  ANDN U17509 ( .A(n17771), .B(n17667), .Z(n17770) );
  XNOR U17510 ( .A(n17769), .B(n17772), .Z(n17667) );
  XNOR U17511 ( .A(n17769), .B(n17665), .Z(n17771) );
  XOR U17512 ( .A(n17773), .B(n17774), .Z(n17665) );
  IV U17513 ( .A(n17775), .Z(n17774) );
  XOR U17514 ( .A(n17776), .B(n17777), .Z(n17769) );
  NANDN U17515 ( .B(n17671), .A(n17778), .Z(n17776) );
  XOR U17516 ( .A(n17777), .B(n17669), .Z(n17778) );
  XOR U17517 ( .A(n17779), .B(n17780), .Z(n17669) );
  IV U17518 ( .A(n17781), .Z(n17780) );
  XNOR U17519 ( .A(n17782), .B(n17777), .Z(n17671) );
  OR U17520 ( .A(n12085), .B(n12086), .Z(n17777) );
  XOR U17521 ( .A(n17783), .B(n17784), .Z(n12085) );
  IV U17522 ( .A(n17785), .Z(n17784) );
  NAND U17523 ( .A(n16747), .B(n17688), .Z(n17782) );
  XOR U17524 ( .A(n16680), .B(n17786), .Z(n16674) );
  IV U17525 ( .A(n16679), .Z(n17786) );
  XNOR U17526 ( .A(n16676), .B(n17276), .Z(n16679) );
  AND U17527 ( .A(n17814), .B(n15896), .Z(n17276) );
  XOR U17528 ( .A(n17787), .B(n17788), .Z(n16676) );
  ANDN U17529 ( .A(n17789), .B(n17678), .Z(n17788) );
  XNOR U17530 ( .A(n17787), .B(n17369), .Z(n17678) );
  AND U17531 ( .A(n17814), .B(n16265), .Z(n17369) );
  XNOR U17532 ( .A(n17787), .B(n17676), .Z(n17789) );
  XOR U17533 ( .A(n17790), .B(n17791), .Z(n17676) );
  IV U17534 ( .A(n17792), .Z(n17791) );
  XOR U17535 ( .A(n17793), .B(n17794), .Z(n17787) );
  ANDN U17536 ( .A(n17795), .B(n17684), .Z(n17794) );
  XNOR U17537 ( .A(n17793), .B(n17472), .Z(n17684) );
  AND U17538 ( .A(n17814), .B(n16657), .Z(n17472) );
  XNOR U17539 ( .A(n17793), .B(n17682), .Z(n17795) );
  XOR U17540 ( .A(n17796), .B(n17797), .Z(n17682) );
  IV U17541 ( .A(n17798), .Z(n17797) );
  XOR U17542 ( .A(n17799), .B(n17800), .Z(n17793) );
  ANDN U17543 ( .A(n17801), .B(n17691), .Z(n17800) );
  XNOR U17544 ( .A(n17799), .B(n17581), .Z(n17691) );
  AND U17545 ( .A(n17814), .B(n17567), .Z(n17581) );
  XNOR U17546 ( .A(n17799), .B(n17689), .Z(n17801) );
  XOR U17547 ( .A(n17802), .B(n17803), .Z(n17689) );
  IV U17548 ( .A(n17804), .Z(n17803) );
  XOR U17549 ( .A(n17805), .B(n17806), .Z(n17799) );
  ANDN U17550 ( .A(n17807), .B(n17698), .Z(n17806) );
  XNOR U17551 ( .A(n17805), .B(n17695), .Z(n17698) );
  AND U17552 ( .A(n17814), .B(n17688), .Z(n17695) );
  XNOR U17553 ( .A(n17805), .B(n17696), .Z(n17807) );
  XOR U17554 ( .A(n17808), .B(n17809), .Z(n17696) );
  IV U17555 ( .A(n17810), .Z(n17809) );
  XOR U17556 ( .A(n17811), .B(n17812), .Z(n17805) );
  ANDN U17557 ( .A(n17813), .B(n17705), .Z(n17812) );
  XNOR U17558 ( .A(n17811), .B(n17814), .Z(n17705) );
  XNOR U17559 ( .A(n17811), .B(n17703), .Z(n17813) );
  XOR U17560 ( .A(n17815), .B(n17816), .Z(n17703) );
  IV U17561 ( .A(n17817), .Z(n17816) );
  XOR U17562 ( .A(n17818), .B(n17819), .Z(n17811) );
  ANDN U17563 ( .A(n17820), .B(n17712), .Z(n17819) );
  XNOR U17564 ( .A(n17818), .B(n17821), .Z(n17712) );
  XNOR U17565 ( .A(n17818), .B(n17710), .Z(n17820) );
  XOR U17566 ( .A(n17822), .B(n17823), .Z(n17710) );
  IV U17567 ( .A(n17824), .Z(n17823) );
  XOR U17568 ( .A(n17825), .B(n17826), .Z(n17818) );
  ANDN U17569 ( .A(n17827), .B(n17719), .Z(n17826) );
  XNOR U17570 ( .A(n17825), .B(n17828), .Z(n17719) );
  XNOR U17571 ( .A(n17825), .B(n17717), .Z(n17827) );
  XOR U17572 ( .A(n17829), .B(n17830), .Z(n17717) );
  IV U17573 ( .A(n17831), .Z(n17830) );
  XOR U17574 ( .A(n17832), .B(n17833), .Z(n17825) );
  ANDN U17575 ( .A(n17834), .B(n17726), .Z(n17833) );
  XNOR U17576 ( .A(n17832), .B(n17835), .Z(n17726) );
  XNOR U17577 ( .A(n17832), .B(n17724), .Z(n17834) );
  XOR U17578 ( .A(n17836), .B(n17837), .Z(n17724) );
  IV U17579 ( .A(n17838), .Z(n17837) );
  XOR U17580 ( .A(n17839), .B(n17840), .Z(n17832) );
  ANDN U17581 ( .A(n17841), .B(n17733), .Z(n17840) );
  XNOR U17582 ( .A(n17839), .B(n17842), .Z(n17733) );
  XNOR U17583 ( .A(n17839), .B(n17731), .Z(n17841) );
  XOR U17584 ( .A(n17843), .B(n17844), .Z(n17731) );
  IV U17585 ( .A(n17845), .Z(n17844) );
  XOR U17586 ( .A(n17846), .B(n17847), .Z(n17839) );
  ANDN U17587 ( .A(n17848), .B(n17740), .Z(n17847) );
  XNOR U17588 ( .A(n17846), .B(n17849), .Z(n17740) );
  XNOR U17589 ( .A(n17846), .B(n17738), .Z(n17848) );
  XOR U17590 ( .A(n17850), .B(n17851), .Z(n17738) );
  IV U17591 ( .A(n17852), .Z(n17851) );
  XOR U17592 ( .A(n17853), .B(n17854), .Z(n17846) );
  ANDN U17593 ( .A(n17855), .B(n17747), .Z(n17854) );
  XNOR U17594 ( .A(n17853), .B(n17856), .Z(n17747) );
  XNOR U17595 ( .A(n17853), .B(n17745), .Z(n17855) );
  XOR U17596 ( .A(n17857), .B(n17858), .Z(n17745) );
  IV U17597 ( .A(n17859), .Z(n17858) );
  XOR U17598 ( .A(n17860), .B(n17861), .Z(n17853) );
  ANDN U17599 ( .A(n17862), .B(n17754), .Z(n17861) );
  XNOR U17600 ( .A(n17860), .B(n17863), .Z(n17754) );
  XNOR U17601 ( .A(n17860), .B(n17752), .Z(n17862) );
  XOR U17602 ( .A(n17864), .B(n17865), .Z(n17752) );
  IV U17603 ( .A(n17866), .Z(n17865) );
  XOR U17604 ( .A(n17867), .B(n17868), .Z(n17860) );
  ANDN U17605 ( .A(n17869), .B(n17761), .Z(n17868) );
  XNOR U17606 ( .A(n17867), .B(n17870), .Z(n17761) );
  XNOR U17607 ( .A(n17867), .B(n17759), .Z(n17869) );
  XOR U17608 ( .A(n17871), .B(n17872), .Z(n17759) );
  IV U17609 ( .A(n17873), .Z(n17872) );
  XOR U17610 ( .A(n17874), .B(n17875), .Z(n17867) );
  ANDN U17611 ( .A(n17876), .B(n17768), .Z(n17875) );
  XNOR U17612 ( .A(n17874), .B(n17877), .Z(n17768) );
  XNOR U17613 ( .A(n17874), .B(n17766), .Z(n17876) );
  XOR U17614 ( .A(n17878), .B(n17879), .Z(n17766) );
  IV U17615 ( .A(n17880), .Z(n17879) );
  XOR U17616 ( .A(n17881), .B(n17882), .Z(n17874) );
  ANDN U17617 ( .A(n17883), .B(n17775), .Z(n17882) );
  XNOR U17618 ( .A(n17881), .B(n17884), .Z(n17775) );
  XNOR U17619 ( .A(n17881), .B(n17773), .Z(n17883) );
  XOR U17620 ( .A(n17885), .B(n17886), .Z(n17773) );
  IV U17621 ( .A(n17887), .Z(n17886) );
  XOR U17622 ( .A(n17888), .B(n17889), .Z(n17881) );
  ANDN U17623 ( .A(n17890), .B(n17781), .Z(n17889) );
  XNOR U17624 ( .A(n17888), .B(n17891), .Z(n17781) );
  XNOR U17625 ( .A(n17888), .B(n17779), .Z(n17890) );
  XOR U17626 ( .A(n17892), .B(n17893), .Z(n17779) );
  IV U17627 ( .A(n17894), .Z(n17893) );
  XOR U17628 ( .A(n17895), .B(n17896), .Z(n17888) );
  NANDN U17629 ( .B(n17785), .A(n17897), .Z(n17895) );
  XOR U17630 ( .A(n17896), .B(n17783), .Z(n17897) );
  XOR U17631 ( .A(n17898), .B(n17899), .Z(n17783) );
  IV U17632 ( .A(n17900), .Z(n17899) );
  XNOR U17633 ( .A(n17901), .B(n17896), .Z(n17785) );
  OR U17634 ( .A(n12218), .B(n12219), .Z(n17896) );
  XOR U17635 ( .A(n17902), .B(n17903), .Z(n12218) );
  IV U17636 ( .A(n17904), .Z(n17903) );
  NAND U17637 ( .A(n16747), .B(n17814), .Z(n17901) );
  XOR U17638 ( .A(n16686), .B(n17905), .Z(n16680) );
  IV U17639 ( .A(n16685), .Z(n17905) );
  XNOR U17640 ( .A(n16682), .B(n17194), .Z(n16685) );
  AND U17641 ( .A(n17945), .B(n15553), .Z(n17194) );
  XOR U17642 ( .A(n17906), .B(n17907), .Z(n16682) );
  ANDN U17643 ( .A(n17908), .B(n17792), .Z(n17907) );
  XNOR U17644 ( .A(n17906), .B(n17280), .Z(n17792) );
  AND U17645 ( .A(n17945), .B(n15896), .Z(n17280) );
  XNOR U17646 ( .A(n17906), .B(n17790), .Z(n17908) );
  XOR U17647 ( .A(n17909), .B(n17910), .Z(n17790) );
  IV U17648 ( .A(n17911), .Z(n17910) );
  XOR U17649 ( .A(n17912), .B(n17913), .Z(n17906) );
  ANDN U17650 ( .A(n17914), .B(n17798), .Z(n17913) );
  XNOR U17651 ( .A(n17912), .B(n17376), .Z(n17798) );
  AND U17652 ( .A(n17945), .B(n16265), .Z(n17376) );
  XNOR U17653 ( .A(n17912), .B(n17796), .Z(n17914) );
  XOR U17654 ( .A(n17915), .B(n17916), .Z(n17796) );
  IV U17655 ( .A(n17917), .Z(n17916) );
  XOR U17656 ( .A(n17918), .B(n17919), .Z(n17912) );
  ANDN U17657 ( .A(n17920), .B(n17804), .Z(n17919) );
  XNOR U17658 ( .A(n17918), .B(n17479), .Z(n17804) );
  AND U17659 ( .A(n17945), .B(n16657), .Z(n17479) );
  XNOR U17660 ( .A(n17918), .B(n17802), .Z(n17920) );
  XOR U17661 ( .A(n17921), .B(n17922), .Z(n17802) );
  IV U17662 ( .A(n17923), .Z(n17922) );
  XOR U17663 ( .A(n17924), .B(n17925), .Z(n17918) );
  ANDN U17664 ( .A(n17926), .B(n17810), .Z(n17925) );
  XNOR U17665 ( .A(n17924), .B(n17588), .Z(n17810) );
  AND U17666 ( .A(n17945), .B(n17567), .Z(n17588) );
  XNOR U17667 ( .A(n17924), .B(n17808), .Z(n17926) );
  XOR U17668 ( .A(n17927), .B(n17928), .Z(n17808) );
  IV U17669 ( .A(n17929), .Z(n17928) );
  XOR U17670 ( .A(n17930), .B(n17931), .Z(n17924) );
  ANDN U17671 ( .A(n17932), .B(n17817), .Z(n17931) );
  XNOR U17672 ( .A(n17930), .B(n17702), .Z(n17817) );
  AND U17673 ( .A(n17945), .B(n17688), .Z(n17702) );
  XNOR U17674 ( .A(n17930), .B(n17815), .Z(n17932) );
  XOR U17675 ( .A(n17933), .B(n17934), .Z(n17815) );
  IV U17676 ( .A(n17935), .Z(n17934) );
  XOR U17677 ( .A(n17936), .B(n17937), .Z(n17930) );
  ANDN U17678 ( .A(n17938), .B(n17824), .Z(n17937) );
  XNOR U17679 ( .A(n17936), .B(n17821), .Z(n17824) );
  AND U17680 ( .A(n17945), .B(n17814), .Z(n17821) );
  XNOR U17681 ( .A(n17936), .B(n17822), .Z(n17938) );
  XOR U17682 ( .A(n17939), .B(n17940), .Z(n17822) );
  IV U17683 ( .A(n17941), .Z(n17940) );
  XOR U17684 ( .A(n17942), .B(n17943), .Z(n17936) );
  ANDN U17685 ( .A(n17944), .B(n17831), .Z(n17943) );
  XNOR U17686 ( .A(n17942), .B(n17945), .Z(n17831) );
  XNOR U17687 ( .A(n17942), .B(n17829), .Z(n17944) );
  XOR U17688 ( .A(n17946), .B(n17947), .Z(n17829) );
  IV U17689 ( .A(n17948), .Z(n17947) );
  XOR U17690 ( .A(n17949), .B(n17950), .Z(n17942) );
  ANDN U17691 ( .A(n17951), .B(n17838), .Z(n17950) );
  XNOR U17692 ( .A(n17949), .B(n17952), .Z(n17838) );
  XNOR U17693 ( .A(n17949), .B(n17836), .Z(n17951) );
  XOR U17694 ( .A(n17953), .B(n17954), .Z(n17836) );
  IV U17695 ( .A(n17955), .Z(n17954) );
  XOR U17696 ( .A(n17956), .B(n17957), .Z(n17949) );
  ANDN U17697 ( .A(n17958), .B(n17845), .Z(n17957) );
  XNOR U17698 ( .A(n17956), .B(n17959), .Z(n17845) );
  XNOR U17699 ( .A(n17956), .B(n17843), .Z(n17958) );
  XOR U17700 ( .A(n17960), .B(n17961), .Z(n17843) );
  IV U17701 ( .A(n17962), .Z(n17961) );
  XOR U17702 ( .A(n17963), .B(n17964), .Z(n17956) );
  ANDN U17703 ( .A(n17965), .B(n17852), .Z(n17964) );
  XNOR U17704 ( .A(n17963), .B(n17966), .Z(n17852) );
  XNOR U17705 ( .A(n17963), .B(n17850), .Z(n17965) );
  XOR U17706 ( .A(n17967), .B(n17968), .Z(n17850) );
  IV U17707 ( .A(n17969), .Z(n17968) );
  XOR U17708 ( .A(n17970), .B(n17971), .Z(n17963) );
  ANDN U17709 ( .A(n17972), .B(n17859), .Z(n17971) );
  XNOR U17710 ( .A(n17970), .B(n17973), .Z(n17859) );
  XNOR U17711 ( .A(n17970), .B(n17857), .Z(n17972) );
  XOR U17712 ( .A(n17974), .B(n17975), .Z(n17857) );
  IV U17713 ( .A(n17976), .Z(n17975) );
  XOR U17714 ( .A(n17977), .B(n17978), .Z(n17970) );
  ANDN U17715 ( .A(n17979), .B(n17866), .Z(n17978) );
  XNOR U17716 ( .A(n17977), .B(n17980), .Z(n17866) );
  XNOR U17717 ( .A(n17977), .B(n17864), .Z(n17979) );
  XOR U17718 ( .A(n17981), .B(n17982), .Z(n17864) );
  IV U17719 ( .A(n17983), .Z(n17982) );
  XOR U17720 ( .A(n17984), .B(n17985), .Z(n17977) );
  ANDN U17721 ( .A(n17986), .B(n17873), .Z(n17985) );
  XNOR U17722 ( .A(n17984), .B(n17987), .Z(n17873) );
  XNOR U17723 ( .A(n17984), .B(n17871), .Z(n17986) );
  XOR U17724 ( .A(n17988), .B(n17989), .Z(n17871) );
  IV U17725 ( .A(n17990), .Z(n17989) );
  XOR U17726 ( .A(n17991), .B(n17992), .Z(n17984) );
  ANDN U17727 ( .A(n17993), .B(n17880), .Z(n17992) );
  XNOR U17728 ( .A(n17991), .B(n17994), .Z(n17880) );
  XNOR U17729 ( .A(n17991), .B(n17878), .Z(n17993) );
  XOR U17730 ( .A(n17995), .B(n17996), .Z(n17878) );
  IV U17731 ( .A(n17997), .Z(n17996) );
  XOR U17732 ( .A(n17998), .B(n17999), .Z(n17991) );
  ANDN U17733 ( .A(n18000), .B(n17887), .Z(n17999) );
  XNOR U17734 ( .A(n17998), .B(n18001), .Z(n17887) );
  XNOR U17735 ( .A(n17998), .B(n17885), .Z(n18000) );
  XOR U17736 ( .A(n18002), .B(n18003), .Z(n17885) );
  IV U17737 ( .A(n18004), .Z(n18003) );
  XOR U17738 ( .A(n18005), .B(n18006), .Z(n17998) );
  ANDN U17739 ( .A(n18007), .B(n17894), .Z(n18006) );
  XNOR U17740 ( .A(n18005), .B(n18008), .Z(n17894) );
  XNOR U17741 ( .A(n18005), .B(n17892), .Z(n18007) );
  XOR U17742 ( .A(n18009), .B(n18010), .Z(n17892) );
  IV U17743 ( .A(n18011), .Z(n18010) );
  XOR U17744 ( .A(n18012), .B(n18013), .Z(n18005) );
  ANDN U17745 ( .A(n18014), .B(n17900), .Z(n18013) );
  XNOR U17746 ( .A(n18012), .B(n18015), .Z(n17900) );
  XNOR U17747 ( .A(n18012), .B(n17898), .Z(n18014) );
  XOR U17748 ( .A(n18016), .B(n18017), .Z(n17898) );
  IV U17749 ( .A(n18018), .Z(n18017) );
  XOR U17750 ( .A(n18019), .B(n18020), .Z(n18012) );
  NANDN U17751 ( .B(n17904), .A(n18021), .Z(n18019) );
  XOR U17752 ( .A(n18020), .B(n17902), .Z(n18021) );
  XOR U17753 ( .A(n18022), .B(n18023), .Z(n17902) );
  IV U17754 ( .A(n18024), .Z(n18023) );
  XNOR U17755 ( .A(n18025), .B(n18020), .Z(n17904) );
  OR U17756 ( .A(n12351), .B(n12352), .Z(n18020) );
  XOR U17757 ( .A(n18026), .B(n18027), .Z(n12351) );
  IV U17758 ( .A(n18028), .Z(n18027) );
  NAND U17759 ( .A(n16747), .B(n17945), .Z(n18025) );
  XOR U17760 ( .A(n16692), .B(n18029), .Z(n16686) );
  IV U17761 ( .A(n16691), .Z(n18029) );
  XNOR U17762 ( .A(n16688), .B(n17119), .Z(n16691) );
  AND U17763 ( .A(n18081), .B(n15236), .Z(n17119) );
  XOR U17764 ( .A(n18030), .B(n18031), .Z(n16688) );
  ANDN U17765 ( .A(n18032), .B(n17911), .Z(n18031) );
  XNOR U17766 ( .A(n18030), .B(n17198), .Z(n17911) );
  AND U17767 ( .A(n18081), .B(n15553), .Z(n17198) );
  XNOR U17768 ( .A(n18030), .B(n17909), .Z(n18032) );
  XOR U17769 ( .A(n18033), .B(n18034), .Z(n17909) );
  IV U17770 ( .A(n18035), .Z(n18034) );
  XOR U17771 ( .A(n18036), .B(n18037), .Z(n18030) );
  ANDN U17772 ( .A(n18038), .B(n17917), .Z(n18037) );
  XNOR U17773 ( .A(n18036), .B(n17287), .Z(n17917) );
  AND U17774 ( .A(n18081), .B(n15896), .Z(n17287) );
  XNOR U17775 ( .A(n18036), .B(n17915), .Z(n18038) );
  XOR U17776 ( .A(n18039), .B(n18040), .Z(n17915) );
  IV U17777 ( .A(n18041), .Z(n18040) );
  XOR U17778 ( .A(n18042), .B(n18043), .Z(n18036) );
  ANDN U17779 ( .A(n18044), .B(n17923), .Z(n18043) );
  XNOR U17780 ( .A(n18042), .B(n17383), .Z(n17923) );
  AND U17781 ( .A(n18081), .B(n16265), .Z(n17383) );
  XNOR U17782 ( .A(n18042), .B(n17921), .Z(n18044) );
  XOR U17783 ( .A(n18045), .B(n18046), .Z(n17921) );
  IV U17784 ( .A(n18047), .Z(n18046) );
  XOR U17785 ( .A(n18048), .B(n18049), .Z(n18042) );
  ANDN U17786 ( .A(n18050), .B(n17929), .Z(n18049) );
  XNOR U17787 ( .A(n18048), .B(n17486), .Z(n17929) );
  AND U17788 ( .A(n18081), .B(n16657), .Z(n17486) );
  XNOR U17789 ( .A(n18048), .B(n17927), .Z(n18050) );
  XOR U17790 ( .A(n18051), .B(n18052), .Z(n17927) );
  IV U17791 ( .A(n18053), .Z(n18052) );
  XOR U17792 ( .A(n18054), .B(n18055), .Z(n18048) );
  ANDN U17793 ( .A(n18056), .B(n17935), .Z(n18055) );
  XNOR U17794 ( .A(n18054), .B(n17595), .Z(n17935) );
  AND U17795 ( .A(n18081), .B(n17567), .Z(n17595) );
  XNOR U17796 ( .A(n18054), .B(n17933), .Z(n18056) );
  XOR U17797 ( .A(n18057), .B(n18058), .Z(n17933) );
  IV U17798 ( .A(n18059), .Z(n18058) );
  XOR U17799 ( .A(n18060), .B(n18061), .Z(n18054) );
  ANDN U17800 ( .A(n18062), .B(n17941), .Z(n18061) );
  XNOR U17801 ( .A(n18060), .B(n17709), .Z(n17941) );
  AND U17802 ( .A(n18081), .B(n17688), .Z(n17709) );
  XNOR U17803 ( .A(n18060), .B(n17939), .Z(n18062) );
  XOR U17804 ( .A(n18063), .B(n18064), .Z(n17939) );
  IV U17805 ( .A(n18065), .Z(n18064) );
  XOR U17806 ( .A(n18066), .B(n18067), .Z(n18060) );
  ANDN U17807 ( .A(n18068), .B(n17948), .Z(n18067) );
  XNOR U17808 ( .A(n18066), .B(n17828), .Z(n17948) );
  AND U17809 ( .A(n18081), .B(n17814), .Z(n17828) );
  XNOR U17810 ( .A(n18066), .B(n17946), .Z(n18068) );
  XOR U17811 ( .A(n18069), .B(n18070), .Z(n17946) );
  IV U17812 ( .A(n18071), .Z(n18070) );
  XOR U17813 ( .A(n18072), .B(n18073), .Z(n18066) );
  ANDN U17814 ( .A(n18074), .B(n17955), .Z(n18073) );
  XNOR U17815 ( .A(n18072), .B(n17952), .Z(n17955) );
  AND U17816 ( .A(n18081), .B(n17945), .Z(n17952) );
  XNOR U17817 ( .A(n18072), .B(n17953), .Z(n18074) );
  XOR U17818 ( .A(n18075), .B(n18076), .Z(n17953) );
  IV U17819 ( .A(n18077), .Z(n18076) );
  XOR U17820 ( .A(n18078), .B(n18079), .Z(n18072) );
  ANDN U17821 ( .A(n18080), .B(n17962), .Z(n18079) );
  XNOR U17822 ( .A(n18078), .B(n18081), .Z(n17962) );
  XNOR U17823 ( .A(n18078), .B(n17960), .Z(n18080) );
  XOR U17824 ( .A(n18082), .B(n18083), .Z(n17960) );
  IV U17825 ( .A(n18084), .Z(n18083) );
  XOR U17826 ( .A(n18085), .B(n18086), .Z(n18078) );
  ANDN U17827 ( .A(n18087), .B(n17969), .Z(n18086) );
  XNOR U17828 ( .A(n18085), .B(n18088), .Z(n17969) );
  XNOR U17829 ( .A(n18085), .B(n17967), .Z(n18087) );
  XOR U17830 ( .A(n18089), .B(n18090), .Z(n17967) );
  IV U17831 ( .A(n18091), .Z(n18090) );
  XOR U17832 ( .A(n18092), .B(n18093), .Z(n18085) );
  ANDN U17833 ( .A(n18094), .B(n17976), .Z(n18093) );
  XNOR U17834 ( .A(n18092), .B(n18095), .Z(n17976) );
  XNOR U17835 ( .A(n18092), .B(n17974), .Z(n18094) );
  XOR U17836 ( .A(n18096), .B(n18097), .Z(n17974) );
  IV U17837 ( .A(n18098), .Z(n18097) );
  XOR U17838 ( .A(n18099), .B(n18100), .Z(n18092) );
  ANDN U17839 ( .A(n18101), .B(n17983), .Z(n18100) );
  XNOR U17840 ( .A(n18099), .B(n18102), .Z(n17983) );
  XNOR U17841 ( .A(n18099), .B(n17981), .Z(n18101) );
  XOR U17842 ( .A(n18103), .B(n18104), .Z(n17981) );
  IV U17843 ( .A(n18105), .Z(n18104) );
  XOR U17844 ( .A(n18106), .B(n18107), .Z(n18099) );
  ANDN U17845 ( .A(n18108), .B(n17990), .Z(n18107) );
  XNOR U17846 ( .A(n18106), .B(n18109), .Z(n17990) );
  XNOR U17847 ( .A(n18106), .B(n17988), .Z(n18108) );
  XOR U17848 ( .A(n18110), .B(n18111), .Z(n17988) );
  IV U17849 ( .A(n18112), .Z(n18111) );
  XOR U17850 ( .A(n18113), .B(n18114), .Z(n18106) );
  ANDN U17851 ( .A(n18115), .B(n17997), .Z(n18114) );
  XNOR U17852 ( .A(n18113), .B(n18116), .Z(n17997) );
  XNOR U17853 ( .A(n18113), .B(n17995), .Z(n18115) );
  XOR U17854 ( .A(n18117), .B(n18118), .Z(n17995) );
  IV U17855 ( .A(n18119), .Z(n18118) );
  XOR U17856 ( .A(n18120), .B(n18121), .Z(n18113) );
  ANDN U17857 ( .A(n18122), .B(n18004), .Z(n18121) );
  XNOR U17858 ( .A(n18120), .B(n18123), .Z(n18004) );
  XNOR U17859 ( .A(n18120), .B(n18002), .Z(n18122) );
  XOR U17860 ( .A(n18124), .B(n18125), .Z(n18002) );
  IV U17861 ( .A(n18126), .Z(n18125) );
  XOR U17862 ( .A(n18127), .B(n18128), .Z(n18120) );
  ANDN U17863 ( .A(n18129), .B(n18011), .Z(n18128) );
  XNOR U17864 ( .A(n18127), .B(n18130), .Z(n18011) );
  XNOR U17865 ( .A(n18127), .B(n18009), .Z(n18129) );
  XOR U17866 ( .A(n18131), .B(n18132), .Z(n18009) );
  IV U17867 ( .A(n18133), .Z(n18132) );
  XOR U17868 ( .A(n18134), .B(n18135), .Z(n18127) );
  ANDN U17869 ( .A(n18136), .B(n18018), .Z(n18135) );
  XNOR U17870 ( .A(n18134), .B(n18137), .Z(n18018) );
  XNOR U17871 ( .A(n18134), .B(n18016), .Z(n18136) );
  XOR U17872 ( .A(n18138), .B(n18139), .Z(n18016) );
  IV U17873 ( .A(n18140), .Z(n18139) );
  XOR U17874 ( .A(n18141), .B(n18142), .Z(n18134) );
  ANDN U17875 ( .A(n18143), .B(n18024), .Z(n18142) );
  XNOR U17876 ( .A(n18141), .B(n18144), .Z(n18024) );
  XNOR U17877 ( .A(n18141), .B(n18022), .Z(n18143) );
  XOR U17878 ( .A(n18145), .B(n18146), .Z(n18022) );
  IV U17879 ( .A(n18147), .Z(n18146) );
  XOR U17880 ( .A(n18148), .B(n18149), .Z(n18141) );
  NANDN U17881 ( .B(n18028), .A(n18150), .Z(n18148) );
  XOR U17882 ( .A(n18149), .B(n18026), .Z(n18150) );
  XOR U17883 ( .A(n18151), .B(n18152), .Z(n18026) );
  IV U17884 ( .A(n18153), .Z(n18152) );
  XNOR U17885 ( .A(n18154), .B(n18149), .Z(n18028) );
  OR U17886 ( .A(n12484), .B(n12485), .Z(n18149) );
  XOR U17887 ( .A(n18155), .B(n18156), .Z(n12484) );
  IV U17888 ( .A(n18157), .Z(n18156) );
  NAND U17889 ( .A(n16747), .B(n18081), .Z(n18154) );
  XOR U17890 ( .A(n16698), .B(n18158), .Z(n16692) );
  IV U17891 ( .A(n16697), .Z(n18158) );
  XNOR U17892 ( .A(n16694), .B(n17051), .Z(n16697) );
  AND U17893 ( .A(n18222), .B(n14945), .Z(n17051) );
  XOR U17894 ( .A(n18159), .B(n18160), .Z(n16694) );
  ANDN U17895 ( .A(n18161), .B(n18035), .Z(n18160) );
  XNOR U17896 ( .A(n18159), .B(n17123), .Z(n18035) );
  AND U17897 ( .A(n18222), .B(n15236), .Z(n17123) );
  XNOR U17898 ( .A(n18159), .B(n18033), .Z(n18161) );
  XOR U17899 ( .A(n18162), .B(n18163), .Z(n18033) );
  IV U17900 ( .A(n18164), .Z(n18163) );
  XOR U17901 ( .A(n18165), .B(n18166), .Z(n18159) );
  ANDN U17902 ( .A(n18167), .B(n18041), .Z(n18166) );
  XNOR U17903 ( .A(n18165), .B(n17205), .Z(n18041) );
  AND U17904 ( .A(n18222), .B(n15553), .Z(n17205) );
  XNOR U17905 ( .A(n18165), .B(n18039), .Z(n18167) );
  XOR U17906 ( .A(n18168), .B(n18169), .Z(n18039) );
  IV U17907 ( .A(n18170), .Z(n18169) );
  XOR U17908 ( .A(n18171), .B(n18172), .Z(n18165) );
  ANDN U17909 ( .A(n18173), .B(n18047), .Z(n18172) );
  XNOR U17910 ( .A(n18171), .B(n17294), .Z(n18047) );
  AND U17911 ( .A(n18222), .B(n15896), .Z(n17294) );
  XNOR U17912 ( .A(n18171), .B(n18045), .Z(n18173) );
  XOR U17913 ( .A(n18174), .B(n18175), .Z(n18045) );
  IV U17914 ( .A(n18176), .Z(n18175) );
  XOR U17915 ( .A(n18177), .B(n18178), .Z(n18171) );
  ANDN U17916 ( .A(n18179), .B(n18053), .Z(n18178) );
  XNOR U17917 ( .A(n18177), .B(n17390), .Z(n18053) );
  AND U17918 ( .A(n18222), .B(n16265), .Z(n17390) );
  XNOR U17919 ( .A(n18177), .B(n18051), .Z(n18179) );
  XOR U17920 ( .A(n18180), .B(n18181), .Z(n18051) );
  IV U17921 ( .A(n18182), .Z(n18181) );
  XOR U17922 ( .A(n18183), .B(n18184), .Z(n18177) );
  ANDN U17923 ( .A(n18185), .B(n18059), .Z(n18184) );
  XNOR U17924 ( .A(n18183), .B(n17493), .Z(n18059) );
  AND U17925 ( .A(n18222), .B(n16657), .Z(n17493) );
  XNOR U17926 ( .A(n18183), .B(n18057), .Z(n18185) );
  XOR U17927 ( .A(n18186), .B(n18187), .Z(n18057) );
  IV U17928 ( .A(n18188), .Z(n18187) );
  XOR U17929 ( .A(n18189), .B(n18190), .Z(n18183) );
  ANDN U17930 ( .A(n18191), .B(n18065), .Z(n18190) );
  XNOR U17931 ( .A(n18189), .B(n17602), .Z(n18065) );
  AND U17932 ( .A(n18222), .B(n17567), .Z(n17602) );
  XNOR U17933 ( .A(n18189), .B(n18063), .Z(n18191) );
  XOR U17934 ( .A(n18192), .B(n18193), .Z(n18063) );
  IV U17935 ( .A(n18194), .Z(n18193) );
  XOR U17936 ( .A(n18195), .B(n18196), .Z(n18189) );
  ANDN U17937 ( .A(n18197), .B(n18071), .Z(n18196) );
  XNOR U17938 ( .A(n18195), .B(n17716), .Z(n18071) );
  AND U17939 ( .A(n18222), .B(n17688), .Z(n17716) );
  XNOR U17940 ( .A(n18195), .B(n18069), .Z(n18197) );
  XOR U17941 ( .A(n18198), .B(n18199), .Z(n18069) );
  IV U17942 ( .A(n18200), .Z(n18199) );
  XOR U17943 ( .A(n18201), .B(n18202), .Z(n18195) );
  ANDN U17944 ( .A(n18203), .B(n18077), .Z(n18202) );
  XNOR U17945 ( .A(n18201), .B(n17835), .Z(n18077) );
  AND U17946 ( .A(n18222), .B(n17814), .Z(n17835) );
  XNOR U17947 ( .A(n18201), .B(n18075), .Z(n18203) );
  XOR U17948 ( .A(n18204), .B(n18205), .Z(n18075) );
  IV U17949 ( .A(n18206), .Z(n18205) );
  XOR U17950 ( .A(n18207), .B(n18208), .Z(n18201) );
  ANDN U17951 ( .A(n18209), .B(n18084), .Z(n18208) );
  XNOR U17952 ( .A(n18207), .B(n17959), .Z(n18084) );
  AND U17953 ( .A(n18222), .B(n17945), .Z(n17959) );
  XNOR U17954 ( .A(n18207), .B(n18082), .Z(n18209) );
  XOR U17955 ( .A(n18210), .B(n18211), .Z(n18082) );
  IV U17956 ( .A(n18212), .Z(n18211) );
  XOR U17957 ( .A(n18213), .B(n18214), .Z(n18207) );
  ANDN U17958 ( .A(n18215), .B(n18091), .Z(n18214) );
  XNOR U17959 ( .A(n18213), .B(n18088), .Z(n18091) );
  AND U17960 ( .A(n18222), .B(n18081), .Z(n18088) );
  XNOR U17961 ( .A(n18213), .B(n18089), .Z(n18215) );
  XOR U17962 ( .A(n18216), .B(n18217), .Z(n18089) );
  IV U17963 ( .A(n18218), .Z(n18217) );
  XOR U17964 ( .A(n18219), .B(n18220), .Z(n18213) );
  ANDN U17965 ( .A(n18221), .B(n18098), .Z(n18220) );
  XNOR U17966 ( .A(n18219), .B(n18222), .Z(n18098) );
  XNOR U17967 ( .A(n18219), .B(n18096), .Z(n18221) );
  XOR U17968 ( .A(n18223), .B(n18224), .Z(n18096) );
  IV U17969 ( .A(n18225), .Z(n18224) );
  XOR U17970 ( .A(n18226), .B(n18227), .Z(n18219) );
  ANDN U17971 ( .A(n18228), .B(n18105), .Z(n18227) );
  XNOR U17972 ( .A(n18226), .B(n18229), .Z(n18105) );
  XNOR U17973 ( .A(n18226), .B(n18103), .Z(n18228) );
  XOR U17974 ( .A(n18230), .B(n18231), .Z(n18103) );
  IV U17975 ( .A(n18232), .Z(n18231) );
  XOR U17976 ( .A(n18233), .B(n18234), .Z(n18226) );
  ANDN U17977 ( .A(n18235), .B(n18112), .Z(n18234) );
  XNOR U17978 ( .A(n18233), .B(n18236), .Z(n18112) );
  XNOR U17979 ( .A(n18233), .B(n18110), .Z(n18235) );
  XOR U17980 ( .A(n18237), .B(n18238), .Z(n18110) );
  IV U17981 ( .A(n18239), .Z(n18238) );
  XOR U17982 ( .A(n18240), .B(n18241), .Z(n18233) );
  ANDN U17983 ( .A(n18242), .B(n18119), .Z(n18241) );
  XNOR U17984 ( .A(n18240), .B(n18243), .Z(n18119) );
  XNOR U17985 ( .A(n18240), .B(n18117), .Z(n18242) );
  XOR U17986 ( .A(n18244), .B(n18245), .Z(n18117) );
  IV U17987 ( .A(n18246), .Z(n18245) );
  XOR U17988 ( .A(n18247), .B(n18248), .Z(n18240) );
  ANDN U17989 ( .A(n18249), .B(n18126), .Z(n18248) );
  XNOR U17990 ( .A(n18247), .B(n18250), .Z(n18126) );
  XNOR U17991 ( .A(n18247), .B(n18124), .Z(n18249) );
  XOR U17992 ( .A(n18251), .B(n18252), .Z(n18124) );
  IV U17993 ( .A(n18253), .Z(n18252) );
  XOR U17994 ( .A(n18254), .B(n18255), .Z(n18247) );
  ANDN U17995 ( .A(n18256), .B(n18133), .Z(n18255) );
  XNOR U17996 ( .A(n18254), .B(n18257), .Z(n18133) );
  XNOR U17997 ( .A(n18254), .B(n18131), .Z(n18256) );
  XOR U17998 ( .A(n18258), .B(n18259), .Z(n18131) );
  IV U17999 ( .A(n18260), .Z(n18259) );
  XOR U18000 ( .A(n18261), .B(n18262), .Z(n18254) );
  ANDN U18001 ( .A(n18263), .B(n18140), .Z(n18262) );
  XNOR U18002 ( .A(n18261), .B(n18264), .Z(n18140) );
  XNOR U18003 ( .A(n18261), .B(n18138), .Z(n18263) );
  XOR U18004 ( .A(n18265), .B(n18266), .Z(n18138) );
  IV U18005 ( .A(n18267), .Z(n18266) );
  XOR U18006 ( .A(n18268), .B(n18269), .Z(n18261) );
  ANDN U18007 ( .A(n18270), .B(n18147), .Z(n18269) );
  XNOR U18008 ( .A(n18268), .B(n18271), .Z(n18147) );
  XNOR U18009 ( .A(n18268), .B(n18145), .Z(n18270) );
  XOR U18010 ( .A(n18272), .B(n18273), .Z(n18145) );
  IV U18011 ( .A(n18274), .Z(n18273) );
  XOR U18012 ( .A(n18275), .B(n18276), .Z(n18268) );
  ANDN U18013 ( .A(n18277), .B(n18153), .Z(n18276) );
  XNOR U18014 ( .A(n18275), .B(n18278), .Z(n18153) );
  XNOR U18015 ( .A(n18275), .B(n18151), .Z(n18277) );
  XOR U18016 ( .A(n18279), .B(n18280), .Z(n18151) );
  IV U18017 ( .A(n18281), .Z(n18280) );
  XOR U18018 ( .A(n18282), .B(n18283), .Z(n18275) );
  NANDN U18019 ( .B(n18157), .A(n18284), .Z(n18282) );
  XOR U18020 ( .A(n18283), .B(n18155), .Z(n18284) );
  XOR U18021 ( .A(n18285), .B(n18286), .Z(n18155) );
  IV U18022 ( .A(n18287), .Z(n18286) );
  XNOR U18023 ( .A(n18288), .B(n18283), .Z(n18157) );
  OR U18024 ( .A(n12615), .B(n12616), .Z(n18283) );
  XOR U18025 ( .A(n18289), .B(n18290), .Z(n12615) );
  IV U18026 ( .A(n18291), .Z(n18290) );
  NAND U18027 ( .A(n16747), .B(n18222), .Z(n18288) );
  XOR U18028 ( .A(n16704), .B(n18292), .Z(n16698) );
  IV U18029 ( .A(n16703), .Z(n18292) );
  XNOR U18030 ( .A(n16700), .B(n16990), .Z(n16703) );
  AND U18031 ( .A(n18368), .B(n14680), .Z(n16990) );
  XOR U18032 ( .A(n18293), .B(n18294), .Z(n16700) );
  ANDN U18033 ( .A(n18295), .B(n18164), .Z(n18294) );
  XNOR U18034 ( .A(n18293), .B(n17055), .Z(n18164) );
  AND U18035 ( .A(n18368), .B(n14945), .Z(n17055) );
  XNOR U18036 ( .A(n18293), .B(n18162), .Z(n18295) );
  XOR U18037 ( .A(n18296), .B(n18297), .Z(n18162) );
  IV U18038 ( .A(n18298), .Z(n18297) );
  XOR U18039 ( .A(n18299), .B(n18300), .Z(n18293) );
  ANDN U18040 ( .A(n18301), .B(n18170), .Z(n18300) );
  XNOR U18041 ( .A(n18299), .B(n17130), .Z(n18170) );
  AND U18042 ( .A(n18368), .B(n15236), .Z(n17130) );
  XNOR U18043 ( .A(n18299), .B(n18168), .Z(n18301) );
  XOR U18044 ( .A(n18302), .B(n18303), .Z(n18168) );
  IV U18045 ( .A(n18304), .Z(n18303) );
  XOR U18046 ( .A(n18305), .B(n18306), .Z(n18299) );
  ANDN U18047 ( .A(n18307), .B(n18176), .Z(n18306) );
  XNOR U18048 ( .A(n18305), .B(n17212), .Z(n18176) );
  AND U18049 ( .A(n18368), .B(n15553), .Z(n17212) );
  XNOR U18050 ( .A(n18305), .B(n18174), .Z(n18307) );
  XOR U18051 ( .A(n18308), .B(n18309), .Z(n18174) );
  IV U18052 ( .A(n18310), .Z(n18309) );
  XOR U18053 ( .A(n18311), .B(n18312), .Z(n18305) );
  ANDN U18054 ( .A(n18313), .B(n18182), .Z(n18312) );
  XNOR U18055 ( .A(n18311), .B(n17301), .Z(n18182) );
  AND U18056 ( .A(n18368), .B(n15896), .Z(n17301) );
  XNOR U18057 ( .A(n18311), .B(n18180), .Z(n18313) );
  XOR U18058 ( .A(n18314), .B(n18315), .Z(n18180) );
  IV U18059 ( .A(n18316), .Z(n18315) );
  XOR U18060 ( .A(n18317), .B(n18318), .Z(n18311) );
  ANDN U18061 ( .A(n18319), .B(n18188), .Z(n18318) );
  XNOR U18062 ( .A(n18317), .B(n17397), .Z(n18188) );
  AND U18063 ( .A(n18368), .B(n16265), .Z(n17397) );
  XNOR U18064 ( .A(n18317), .B(n18186), .Z(n18319) );
  XOR U18065 ( .A(n18320), .B(n18321), .Z(n18186) );
  IV U18066 ( .A(n18322), .Z(n18321) );
  XOR U18067 ( .A(n18323), .B(n18324), .Z(n18317) );
  ANDN U18068 ( .A(n18325), .B(n18194), .Z(n18324) );
  XNOR U18069 ( .A(n18323), .B(n17500), .Z(n18194) );
  AND U18070 ( .A(n18368), .B(n16657), .Z(n17500) );
  XNOR U18071 ( .A(n18323), .B(n18192), .Z(n18325) );
  XOR U18072 ( .A(n18326), .B(n18327), .Z(n18192) );
  IV U18073 ( .A(n18328), .Z(n18327) );
  XOR U18074 ( .A(n18329), .B(n18330), .Z(n18323) );
  ANDN U18075 ( .A(n18331), .B(n18200), .Z(n18330) );
  XNOR U18076 ( .A(n18329), .B(n17609), .Z(n18200) );
  AND U18077 ( .A(n18368), .B(n17567), .Z(n17609) );
  XNOR U18078 ( .A(n18329), .B(n18198), .Z(n18331) );
  XOR U18079 ( .A(n18332), .B(n18333), .Z(n18198) );
  IV U18080 ( .A(n18334), .Z(n18333) );
  XOR U18081 ( .A(n18335), .B(n18336), .Z(n18329) );
  ANDN U18082 ( .A(n18337), .B(n18206), .Z(n18336) );
  XNOR U18083 ( .A(n18335), .B(n17723), .Z(n18206) );
  AND U18084 ( .A(n18368), .B(n17688), .Z(n17723) );
  XNOR U18085 ( .A(n18335), .B(n18204), .Z(n18337) );
  XOR U18086 ( .A(n18338), .B(n18339), .Z(n18204) );
  IV U18087 ( .A(n18340), .Z(n18339) );
  XOR U18088 ( .A(n18341), .B(n18342), .Z(n18335) );
  ANDN U18089 ( .A(n18343), .B(n18212), .Z(n18342) );
  XNOR U18090 ( .A(n18341), .B(n17842), .Z(n18212) );
  AND U18091 ( .A(n18368), .B(n17814), .Z(n17842) );
  XNOR U18092 ( .A(n18341), .B(n18210), .Z(n18343) );
  XOR U18093 ( .A(n18344), .B(n18345), .Z(n18210) );
  IV U18094 ( .A(n18346), .Z(n18345) );
  XOR U18095 ( .A(n18347), .B(n18348), .Z(n18341) );
  ANDN U18096 ( .A(n18349), .B(n18218), .Z(n18348) );
  XNOR U18097 ( .A(n18347), .B(n17966), .Z(n18218) );
  AND U18098 ( .A(n18368), .B(n17945), .Z(n17966) );
  XNOR U18099 ( .A(n18347), .B(n18216), .Z(n18349) );
  XOR U18100 ( .A(n18350), .B(n18351), .Z(n18216) );
  IV U18101 ( .A(n18352), .Z(n18351) );
  XOR U18102 ( .A(n18353), .B(n18354), .Z(n18347) );
  ANDN U18103 ( .A(n18355), .B(n18225), .Z(n18354) );
  XNOR U18104 ( .A(n18353), .B(n18095), .Z(n18225) );
  AND U18105 ( .A(n18368), .B(n18081), .Z(n18095) );
  XNOR U18106 ( .A(n18353), .B(n18223), .Z(n18355) );
  XOR U18107 ( .A(n18356), .B(n18357), .Z(n18223) );
  IV U18108 ( .A(n18358), .Z(n18357) );
  XOR U18109 ( .A(n18359), .B(n18360), .Z(n18353) );
  ANDN U18110 ( .A(n18361), .B(n18232), .Z(n18360) );
  XNOR U18111 ( .A(n18359), .B(n18229), .Z(n18232) );
  AND U18112 ( .A(n18368), .B(n18222), .Z(n18229) );
  XNOR U18113 ( .A(n18359), .B(n18230), .Z(n18361) );
  XOR U18114 ( .A(n18362), .B(n18363), .Z(n18230) );
  IV U18115 ( .A(n18364), .Z(n18363) );
  XOR U18116 ( .A(n18365), .B(n18366), .Z(n18359) );
  ANDN U18117 ( .A(n18367), .B(n18239), .Z(n18366) );
  XNOR U18118 ( .A(n18365), .B(n18368), .Z(n18239) );
  XNOR U18119 ( .A(n18365), .B(n18237), .Z(n18367) );
  XOR U18120 ( .A(n18369), .B(n18370), .Z(n18237) );
  IV U18121 ( .A(n18371), .Z(n18370) );
  XOR U18122 ( .A(n18372), .B(n18373), .Z(n18365) );
  ANDN U18123 ( .A(n18374), .B(n18246), .Z(n18373) );
  XNOR U18124 ( .A(n18372), .B(n18375), .Z(n18246) );
  XNOR U18125 ( .A(n18372), .B(n18244), .Z(n18374) );
  XOR U18126 ( .A(n18376), .B(n18377), .Z(n18244) );
  IV U18127 ( .A(n18378), .Z(n18377) );
  XOR U18128 ( .A(n18379), .B(n18380), .Z(n18372) );
  ANDN U18129 ( .A(n18381), .B(n18253), .Z(n18380) );
  XNOR U18130 ( .A(n18379), .B(n18382), .Z(n18253) );
  XNOR U18131 ( .A(n18379), .B(n18251), .Z(n18381) );
  XOR U18132 ( .A(n18383), .B(n18384), .Z(n18251) );
  IV U18133 ( .A(n18385), .Z(n18384) );
  XOR U18134 ( .A(n18386), .B(n18387), .Z(n18379) );
  ANDN U18135 ( .A(n18388), .B(n18260), .Z(n18387) );
  XNOR U18136 ( .A(n18386), .B(n18389), .Z(n18260) );
  XNOR U18137 ( .A(n18386), .B(n18258), .Z(n18388) );
  XOR U18138 ( .A(n18390), .B(n18391), .Z(n18258) );
  IV U18139 ( .A(n18392), .Z(n18391) );
  XOR U18140 ( .A(n18393), .B(n18394), .Z(n18386) );
  ANDN U18141 ( .A(n18395), .B(n18267), .Z(n18394) );
  XNOR U18142 ( .A(n18393), .B(n18396), .Z(n18267) );
  XNOR U18143 ( .A(n18393), .B(n18265), .Z(n18395) );
  XOR U18144 ( .A(n18397), .B(n18398), .Z(n18265) );
  IV U18145 ( .A(n18399), .Z(n18398) );
  XOR U18146 ( .A(n18400), .B(n18401), .Z(n18393) );
  ANDN U18147 ( .A(n18402), .B(n18274), .Z(n18401) );
  XNOR U18148 ( .A(n18400), .B(n18403), .Z(n18274) );
  XNOR U18149 ( .A(n18400), .B(n18272), .Z(n18402) );
  XOR U18150 ( .A(n18404), .B(n18405), .Z(n18272) );
  IV U18151 ( .A(n18406), .Z(n18405) );
  XOR U18152 ( .A(n18407), .B(n18408), .Z(n18400) );
  ANDN U18153 ( .A(n18409), .B(n18281), .Z(n18408) );
  XNOR U18154 ( .A(n18407), .B(n18410), .Z(n18281) );
  XNOR U18155 ( .A(n18407), .B(n18279), .Z(n18409) );
  XOR U18156 ( .A(n18411), .B(n18412), .Z(n18279) );
  IV U18157 ( .A(n18413), .Z(n18412) );
  XOR U18158 ( .A(n18414), .B(n18415), .Z(n18407) );
  ANDN U18159 ( .A(n18416), .B(n18287), .Z(n18415) );
  XNOR U18160 ( .A(n18414), .B(n18417), .Z(n18287) );
  XNOR U18161 ( .A(n18414), .B(n18285), .Z(n18416) );
  XOR U18162 ( .A(n18418), .B(n18419), .Z(n18285) );
  IV U18163 ( .A(n18420), .Z(n18419) );
  XOR U18164 ( .A(n18421), .B(n18422), .Z(n18414) );
  NANDN U18165 ( .B(n18291), .A(n18423), .Z(n18421) );
  XOR U18166 ( .A(n18422), .B(n18289), .Z(n18423) );
  XOR U18167 ( .A(n18424), .B(n18425), .Z(n18289) );
  IV U18168 ( .A(n18426), .Z(n18425) );
  XNOR U18169 ( .A(n18427), .B(n18422), .Z(n18291) );
  OR U18170 ( .A(n12739), .B(n12740), .Z(n18422) );
  XOR U18171 ( .A(n18428), .B(n18429), .Z(n12739) );
  IV U18172 ( .A(n18430), .Z(n18429) );
  NAND U18173 ( .A(n16747), .B(n18368), .Z(n18427) );
  XOR U18174 ( .A(n16710), .B(n18431), .Z(n16704) );
  IV U18175 ( .A(n16709), .Z(n18431) );
  XNOR U18176 ( .A(n16706), .B(n16936), .Z(n16709) );
  AND U18177 ( .A(n18519), .B(n14441), .Z(n16936) );
  XOR U18178 ( .A(n18432), .B(n18433), .Z(n16706) );
  ANDN U18179 ( .A(n18434), .B(n18298), .Z(n18433) );
  XNOR U18180 ( .A(n18432), .B(n16994), .Z(n18298) );
  AND U18181 ( .A(n18519), .B(n14680), .Z(n16994) );
  XNOR U18182 ( .A(n18432), .B(n18296), .Z(n18434) );
  XOR U18183 ( .A(n18435), .B(n18436), .Z(n18296) );
  IV U18184 ( .A(n18437), .Z(n18436) );
  XOR U18185 ( .A(n18438), .B(n18439), .Z(n18432) );
  ANDN U18186 ( .A(n18440), .B(n18304), .Z(n18439) );
  XNOR U18187 ( .A(n18438), .B(n17062), .Z(n18304) );
  AND U18188 ( .A(n18519), .B(n14945), .Z(n17062) );
  XNOR U18189 ( .A(n18438), .B(n18302), .Z(n18440) );
  XOR U18190 ( .A(n18441), .B(n18442), .Z(n18302) );
  IV U18191 ( .A(n18443), .Z(n18442) );
  XOR U18192 ( .A(n18444), .B(n18445), .Z(n18438) );
  ANDN U18193 ( .A(n18446), .B(n18310), .Z(n18445) );
  XNOR U18194 ( .A(n18444), .B(n17137), .Z(n18310) );
  AND U18195 ( .A(n18519), .B(n15236), .Z(n17137) );
  XNOR U18196 ( .A(n18444), .B(n18308), .Z(n18446) );
  XOR U18197 ( .A(n18447), .B(n18448), .Z(n18308) );
  IV U18198 ( .A(n18449), .Z(n18448) );
  XOR U18199 ( .A(n18450), .B(n18451), .Z(n18444) );
  ANDN U18200 ( .A(n18452), .B(n18316), .Z(n18451) );
  XNOR U18201 ( .A(n18450), .B(n17219), .Z(n18316) );
  AND U18202 ( .A(n18519), .B(n15553), .Z(n17219) );
  XNOR U18203 ( .A(n18450), .B(n18314), .Z(n18452) );
  XOR U18204 ( .A(n18453), .B(n18454), .Z(n18314) );
  IV U18205 ( .A(n18455), .Z(n18454) );
  XOR U18206 ( .A(n18456), .B(n18457), .Z(n18450) );
  ANDN U18207 ( .A(n18458), .B(n18322), .Z(n18457) );
  XNOR U18208 ( .A(n18456), .B(n17308), .Z(n18322) );
  AND U18209 ( .A(n18519), .B(n15896), .Z(n17308) );
  XNOR U18210 ( .A(n18456), .B(n18320), .Z(n18458) );
  XOR U18211 ( .A(n18459), .B(n18460), .Z(n18320) );
  IV U18212 ( .A(n18461), .Z(n18460) );
  XOR U18213 ( .A(n18462), .B(n18463), .Z(n18456) );
  ANDN U18214 ( .A(n18464), .B(n18328), .Z(n18463) );
  XNOR U18215 ( .A(n18462), .B(n17404), .Z(n18328) );
  AND U18216 ( .A(n18519), .B(n16265), .Z(n17404) );
  XNOR U18217 ( .A(n18462), .B(n18326), .Z(n18464) );
  XOR U18218 ( .A(n18465), .B(n18466), .Z(n18326) );
  IV U18219 ( .A(n18467), .Z(n18466) );
  XOR U18220 ( .A(n18468), .B(n18469), .Z(n18462) );
  ANDN U18221 ( .A(n18470), .B(n18334), .Z(n18469) );
  XNOR U18222 ( .A(n18468), .B(n17507), .Z(n18334) );
  AND U18223 ( .A(n18519), .B(n16657), .Z(n17507) );
  XNOR U18224 ( .A(n18468), .B(n18332), .Z(n18470) );
  XOR U18225 ( .A(n18471), .B(n18472), .Z(n18332) );
  IV U18226 ( .A(n18473), .Z(n18472) );
  XOR U18227 ( .A(n18474), .B(n18475), .Z(n18468) );
  ANDN U18228 ( .A(n18476), .B(n18340), .Z(n18475) );
  XNOR U18229 ( .A(n18474), .B(n17616), .Z(n18340) );
  AND U18230 ( .A(n18519), .B(n17567), .Z(n17616) );
  XNOR U18231 ( .A(n18474), .B(n18338), .Z(n18476) );
  XOR U18232 ( .A(n18477), .B(n18478), .Z(n18338) );
  IV U18233 ( .A(n18479), .Z(n18478) );
  XOR U18234 ( .A(n18480), .B(n18481), .Z(n18474) );
  ANDN U18235 ( .A(n18482), .B(n18346), .Z(n18481) );
  XNOR U18236 ( .A(n18480), .B(n17730), .Z(n18346) );
  AND U18237 ( .A(n18519), .B(n17688), .Z(n17730) );
  XNOR U18238 ( .A(n18480), .B(n18344), .Z(n18482) );
  XOR U18239 ( .A(n18483), .B(n18484), .Z(n18344) );
  IV U18240 ( .A(n18485), .Z(n18484) );
  XOR U18241 ( .A(n18486), .B(n18487), .Z(n18480) );
  ANDN U18242 ( .A(n18488), .B(n18352), .Z(n18487) );
  XNOR U18243 ( .A(n18486), .B(n17849), .Z(n18352) );
  AND U18244 ( .A(n18519), .B(n17814), .Z(n17849) );
  XNOR U18245 ( .A(n18486), .B(n18350), .Z(n18488) );
  XOR U18246 ( .A(n18489), .B(n18490), .Z(n18350) );
  IV U18247 ( .A(n18491), .Z(n18490) );
  XOR U18248 ( .A(n18492), .B(n18493), .Z(n18486) );
  ANDN U18249 ( .A(n18494), .B(n18358), .Z(n18493) );
  XNOR U18250 ( .A(n18492), .B(n17973), .Z(n18358) );
  AND U18251 ( .A(n18519), .B(n17945), .Z(n17973) );
  XNOR U18252 ( .A(n18492), .B(n18356), .Z(n18494) );
  XOR U18253 ( .A(n18495), .B(n18496), .Z(n18356) );
  IV U18254 ( .A(n18497), .Z(n18496) );
  XOR U18255 ( .A(n18498), .B(n18499), .Z(n18492) );
  ANDN U18256 ( .A(n18500), .B(n18364), .Z(n18499) );
  XNOR U18257 ( .A(n18498), .B(n18102), .Z(n18364) );
  AND U18258 ( .A(n18519), .B(n18081), .Z(n18102) );
  XNOR U18259 ( .A(n18498), .B(n18362), .Z(n18500) );
  XOR U18260 ( .A(n18501), .B(n18502), .Z(n18362) );
  IV U18261 ( .A(n18503), .Z(n18502) );
  XOR U18262 ( .A(n18504), .B(n18505), .Z(n18498) );
  ANDN U18263 ( .A(n18506), .B(n18371), .Z(n18505) );
  XNOR U18264 ( .A(n18504), .B(n18236), .Z(n18371) );
  AND U18265 ( .A(n18519), .B(n18222), .Z(n18236) );
  XNOR U18266 ( .A(n18504), .B(n18369), .Z(n18506) );
  XOR U18267 ( .A(n18507), .B(n18508), .Z(n18369) );
  IV U18268 ( .A(n18509), .Z(n18508) );
  XOR U18269 ( .A(n18510), .B(n18511), .Z(n18504) );
  ANDN U18270 ( .A(n18512), .B(n18378), .Z(n18511) );
  XNOR U18271 ( .A(n18510), .B(n18375), .Z(n18378) );
  AND U18272 ( .A(n18519), .B(n18368), .Z(n18375) );
  XNOR U18273 ( .A(n18510), .B(n18376), .Z(n18512) );
  XOR U18274 ( .A(n18513), .B(n18514), .Z(n18376) );
  IV U18275 ( .A(n18515), .Z(n18514) );
  XOR U18276 ( .A(n18516), .B(n18517), .Z(n18510) );
  ANDN U18277 ( .A(n18518), .B(n18385), .Z(n18517) );
  XNOR U18278 ( .A(n18516), .B(n18519), .Z(n18385) );
  XNOR U18279 ( .A(n18516), .B(n18383), .Z(n18518) );
  XOR U18280 ( .A(n18520), .B(n18521), .Z(n18383) );
  IV U18281 ( .A(n18522), .Z(n18521) );
  XOR U18282 ( .A(n18523), .B(n18524), .Z(n18516) );
  ANDN U18283 ( .A(n18525), .B(n18392), .Z(n18524) );
  XNOR U18284 ( .A(n18523), .B(n18526), .Z(n18392) );
  XNOR U18285 ( .A(n18523), .B(n18390), .Z(n18525) );
  XOR U18286 ( .A(n18527), .B(n18528), .Z(n18390) );
  IV U18287 ( .A(n18529), .Z(n18528) );
  XOR U18288 ( .A(n18530), .B(n18531), .Z(n18523) );
  ANDN U18289 ( .A(n18532), .B(n18399), .Z(n18531) );
  XNOR U18290 ( .A(n18530), .B(n18533), .Z(n18399) );
  XNOR U18291 ( .A(n18530), .B(n18397), .Z(n18532) );
  XOR U18292 ( .A(n18534), .B(n18535), .Z(n18397) );
  IV U18293 ( .A(n18536), .Z(n18535) );
  XOR U18294 ( .A(n18537), .B(n18538), .Z(n18530) );
  ANDN U18295 ( .A(n18539), .B(n18406), .Z(n18538) );
  XNOR U18296 ( .A(n18537), .B(n18540), .Z(n18406) );
  XNOR U18297 ( .A(n18537), .B(n18404), .Z(n18539) );
  XOR U18298 ( .A(n18541), .B(n18542), .Z(n18404) );
  IV U18299 ( .A(n18543), .Z(n18542) );
  XOR U18300 ( .A(n18544), .B(n18545), .Z(n18537) );
  ANDN U18301 ( .A(n18546), .B(n18413), .Z(n18545) );
  XNOR U18302 ( .A(n18544), .B(n18547), .Z(n18413) );
  XNOR U18303 ( .A(n18544), .B(n18411), .Z(n18546) );
  XOR U18304 ( .A(n18548), .B(n18549), .Z(n18411) );
  IV U18305 ( .A(n18550), .Z(n18549) );
  XOR U18306 ( .A(n18551), .B(n18552), .Z(n18544) );
  ANDN U18307 ( .A(n18553), .B(n18420), .Z(n18552) );
  XNOR U18308 ( .A(n18551), .B(n18554), .Z(n18420) );
  XNOR U18309 ( .A(n18551), .B(n18418), .Z(n18553) );
  XOR U18310 ( .A(n18555), .B(n18556), .Z(n18418) );
  IV U18311 ( .A(n18557), .Z(n18556) );
  XOR U18312 ( .A(n18558), .B(n18559), .Z(n18551) );
  ANDN U18313 ( .A(n18560), .B(n18426), .Z(n18559) );
  XNOR U18314 ( .A(n18558), .B(n18561), .Z(n18426) );
  XNOR U18315 ( .A(n18558), .B(n18424), .Z(n18560) );
  XOR U18316 ( .A(n18562), .B(n18563), .Z(n18424) );
  IV U18317 ( .A(n18564), .Z(n18563) );
  XOR U18318 ( .A(n18565), .B(n18566), .Z(n18558) );
  NANDN U18319 ( .B(n18430), .A(n18567), .Z(n18565) );
  XOR U18320 ( .A(n18566), .B(n18428), .Z(n18567) );
  XOR U18321 ( .A(n18568), .B(n18569), .Z(n18428) );
  IV U18322 ( .A(n18570), .Z(n18569) );
  XNOR U18323 ( .A(n18571), .B(n18566), .Z(n18430) );
  OR U18324 ( .A(n12858), .B(n12859), .Z(n18566) );
  XOR U18325 ( .A(n18572), .B(n18573), .Z(n12858) );
  IV U18326 ( .A(n18574), .Z(n18573) );
  NAND U18327 ( .A(n16747), .B(n18519), .Z(n18571) );
  XOR U18328 ( .A(n16716), .B(n18575), .Z(n16710) );
  IV U18329 ( .A(n16715), .Z(n18575) );
  XNOR U18330 ( .A(n16712), .B(n16889), .Z(n16715) );
  AND U18331 ( .A(n18675), .B(n14228), .Z(n16889) );
  XOR U18332 ( .A(n18576), .B(n18577), .Z(n16712) );
  ANDN U18333 ( .A(n18578), .B(n18437), .Z(n18577) );
  XNOR U18334 ( .A(n18576), .B(n16940), .Z(n18437) );
  AND U18335 ( .A(n18675), .B(n14441), .Z(n16940) );
  XNOR U18336 ( .A(n18576), .B(n18435), .Z(n18578) );
  XOR U18337 ( .A(n18579), .B(n18580), .Z(n18435) );
  IV U18338 ( .A(n18581), .Z(n18580) );
  XOR U18339 ( .A(n18582), .B(n18583), .Z(n18576) );
  ANDN U18340 ( .A(n18584), .B(n18443), .Z(n18583) );
  XNOR U18341 ( .A(n18582), .B(n17001), .Z(n18443) );
  AND U18342 ( .A(n18675), .B(n14680), .Z(n17001) );
  XNOR U18343 ( .A(n18582), .B(n18441), .Z(n18584) );
  XOR U18344 ( .A(n18585), .B(n18586), .Z(n18441) );
  IV U18345 ( .A(n18587), .Z(n18586) );
  XOR U18346 ( .A(n18588), .B(n18589), .Z(n18582) );
  ANDN U18347 ( .A(n18590), .B(n18449), .Z(n18589) );
  XNOR U18348 ( .A(n18588), .B(n17069), .Z(n18449) );
  AND U18349 ( .A(n18675), .B(n14945), .Z(n17069) );
  XNOR U18350 ( .A(n18588), .B(n18447), .Z(n18590) );
  XOR U18351 ( .A(n18591), .B(n18592), .Z(n18447) );
  IV U18352 ( .A(n18593), .Z(n18592) );
  XOR U18353 ( .A(n18594), .B(n18595), .Z(n18588) );
  ANDN U18354 ( .A(n18596), .B(n18455), .Z(n18595) );
  XNOR U18355 ( .A(n18594), .B(n17144), .Z(n18455) );
  AND U18356 ( .A(n18675), .B(n15236), .Z(n17144) );
  XNOR U18357 ( .A(n18594), .B(n18453), .Z(n18596) );
  XOR U18358 ( .A(n18597), .B(n18598), .Z(n18453) );
  IV U18359 ( .A(n18599), .Z(n18598) );
  XOR U18360 ( .A(n18600), .B(n18601), .Z(n18594) );
  ANDN U18361 ( .A(n18602), .B(n18461), .Z(n18601) );
  XNOR U18362 ( .A(n18600), .B(n17226), .Z(n18461) );
  AND U18363 ( .A(n18675), .B(n15553), .Z(n17226) );
  XNOR U18364 ( .A(n18600), .B(n18459), .Z(n18602) );
  XOR U18365 ( .A(n18603), .B(n18604), .Z(n18459) );
  IV U18366 ( .A(n18605), .Z(n18604) );
  XOR U18367 ( .A(n18606), .B(n18607), .Z(n18600) );
  ANDN U18368 ( .A(n18608), .B(n18467), .Z(n18607) );
  XNOR U18369 ( .A(n18606), .B(n17315), .Z(n18467) );
  AND U18370 ( .A(n18675), .B(n15896), .Z(n17315) );
  XNOR U18371 ( .A(n18606), .B(n18465), .Z(n18608) );
  XOR U18372 ( .A(n18609), .B(n18610), .Z(n18465) );
  IV U18373 ( .A(n18611), .Z(n18610) );
  XOR U18374 ( .A(n18612), .B(n18613), .Z(n18606) );
  ANDN U18375 ( .A(n18614), .B(n18473), .Z(n18613) );
  XNOR U18376 ( .A(n18612), .B(n17411), .Z(n18473) );
  AND U18377 ( .A(n18675), .B(n16265), .Z(n17411) );
  XNOR U18378 ( .A(n18612), .B(n18471), .Z(n18614) );
  XOR U18379 ( .A(n18615), .B(n18616), .Z(n18471) );
  IV U18380 ( .A(n18617), .Z(n18616) );
  XOR U18381 ( .A(n18618), .B(n18619), .Z(n18612) );
  ANDN U18382 ( .A(n18620), .B(n18479), .Z(n18619) );
  XNOR U18383 ( .A(n18618), .B(n17514), .Z(n18479) );
  AND U18384 ( .A(n18675), .B(n16657), .Z(n17514) );
  XNOR U18385 ( .A(n18618), .B(n18477), .Z(n18620) );
  XOR U18386 ( .A(n18621), .B(n18622), .Z(n18477) );
  IV U18387 ( .A(n18623), .Z(n18622) );
  XOR U18388 ( .A(n18624), .B(n18625), .Z(n18618) );
  ANDN U18389 ( .A(n18626), .B(n18485), .Z(n18625) );
  XNOR U18390 ( .A(n18624), .B(n17623), .Z(n18485) );
  AND U18391 ( .A(n18675), .B(n17567), .Z(n17623) );
  XNOR U18392 ( .A(n18624), .B(n18483), .Z(n18626) );
  XOR U18393 ( .A(n18627), .B(n18628), .Z(n18483) );
  IV U18394 ( .A(n18629), .Z(n18628) );
  XOR U18395 ( .A(n18630), .B(n18631), .Z(n18624) );
  ANDN U18396 ( .A(n18632), .B(n18491), .Z(n18631) );
  XNOR U18397 ( .A(n18630), .B(n17737), .Z(n18491) );
  AND U18398 ( .A(n18675), .B(n17688), .Z(n17737) );
  XNOR U18399 ( .A(n18630), .B(n18489), .Z(n18632) );
  XOR U18400 ( .A(n18633), .B(n18634), .Z(n18489) );
  IV U18401 ( .A(n18635), .Z(n18634) );
  XOR U18402 ( .A(n18636), .B(n18637), .Z(n18630) );
  ANDN U18403 ( .A(n18638), .B(n18497), .Z(n18637) );
  XNOR U18404 ( .A(n18636), .B(n17856), .Z(n18497) );
  AND U18405 ( .A(n18675), .B(n17814), .Z(n17856) );
  XNOR U18406 ( .A(n18636), .B(n18495), .Z(n18638) );
  XOR U18407 ( .A(n18639), .B(n18640), .Z(n18495) );
  IV U18408 ( .A(n18641), .Z(n18640) );
  XOR U18409 ( .A(n18642), .B(n18643), .Z(n18636) );
  ANDN U18410 ( .A(n18644), .B(n18503), .Z(n18643) );
  XNOR U18411 ( .A(n18642), .B(n17980), .Z(n18503) );
  AND U18412 ( .A(n18675), .B(n17945), .Z(n17980) );
  XNOR U18413 ( .A(n18642), .B(n18501), .Z(n18644) );
  XOR U18414 ( .A(n18645), .B(n18646), .Z(n18501) );
  IV U18415 ( .A(n18647), .Z(n18646) );
  XOR U18416 ( .A(n18648), .B(n18649), .Z(n18642) );
  ANDN U18417 ( .A(n18650), .B(n18509), .Z(n18649) );
  XNOR U18418 ( .A(n18648), .B(n18109), .Z(n18509) );
  AND U18419 ( .A(n18675), .B(n18081), .Z(n18109) );
  XNOR U18420 ( .A(n18648), .B(n18507), .Z(n18650) );
  XOR U18421 ( .A(n18651), .B(n18652), .Z(n18507) );
  IV U18422 ( .A(n18653), .Z(n18652) );
  XOR U18423 ( .A(n18654), .B(n18655), .Z(n18648) );
  ANDN U18424 ( .A(n18656), .B(n18515), .Z(n18655) );
  XNOR U18425 ( .A(n18654), .B(n18243), .Z(n18515) );
  AND U18426 ( .A(n18675), .B(n18222), .Z(n18243) );
  XNOR U18427 ( .A(n18654), .B(n18513), .Z(n18656) );
  XOR U18428 ( .A(n18657), .B(n18658), .Z(n18513) );
  IV U18429 ( .A(n18659), .Z(n18658) );
  XOR U18430 ( .A(n18660), .B(n18661), .Z(n18654) );
  ANDN U18431 ( .A(n18662), .B(n18522), .Z(n18661) );
  XNOR U18432 ( .A(n18660), .B(n18382), .Z(n18522) );
  AND U18433 ( .A(n18675), .B(n18368), .Z(n18382) );
  XNOR U18434 ( .A(n18660), .B(n18520), .Z(n18662) );
  XOR U18435 ( .A(n18663), .B(n18664), .Z(n18520) );
  IV U18436 ( .A(n18665), .Z(n18664) );
  XOR U18437 ( .A(n18666), .B(n18667), .Z(n18660) );
  ANDN U18438 ( .A(n18668), .B(n18529), .Z(n18667) );
  XNOR U18439 ( .A(n18666), .B(n18526), .Z(n18529) );
  AND U18440 ( .A(n18675), .B(n18519), .Z(n18526) );
  XNOR U18441 ( .A(n18666), .B(n18527), .Z(n18668) );
  XOR U18442 ( .A(n18669), .B(n18670), .Z(n18527) );
  IV U18443 ( .A(n18671), .Z(n18670) );
  XOR U18444 ( .A(n18672), .B(n18673), .Z(n18666) );
  ANDN U18445 ( .A(n18674), .B(n18536), .Z(n18673) );
  XNOR U18446 ( .A(n18672), .B(n18675), .Z(n18536) );
  XNOR U18447 ( .A(n18672), .B(n18534), .Z(n18674) );
  XOR U18448 ( .A(n18676), .B(n18677), .Z(n18534) );
  IV U18449 ( .A(n18678), .Z(n18677) );
  XOR U18450 ( .A(n18679), .B(n18680), .Z(n18672) );
  ANDN U18451 ( .A(n18681), .B(n18543), .Z(n18680) );
  XNOR U18452 ( .A(n18679), .B(n18682), .Z(n18543) );
  XNOR U18453 ( .A(n18679), .B(n18541), .Z(n18681) );
  XOR U18454 ( .A(n18683), .B(n18684), .Z(n18541) );
  IV U18455 ( .A(n18685), .Z(n18684) );
  XOR U18456 ( .A(n18686), .B(n18687), .Z(n18679) );
  ANDN U18457 ( .A(n18688), .B(n18550), .Z(n18687) );
  XNOR U18458 ( .A(n18686), .B(n18689), .Z(n18550) );
  XNOR U18459 ( .A(n18686), .B(n18548), .Z(n18688) );
  XOR U18460 ( .A(n18690), .B(n18691), .Z(n18548) );
  IV U18461 ( .A(n18692), .Z(n18691) );
  XOR U18462 ( .A(n18693), .B(n18694), .Z(n18686) );
  ANDN U18463 ( .A(n18695), .B(n18557), .Z(n18694) );
  XNOR U18464 ( .A(n18693), .B(n18696), .Z(n18557) );
  XNOR U18465 ( .A(n18693), .B(n18555), .Z(n18695) );
  XOR U18466 ( .A(n18697), .B(n18698), .Z(n18555) );
  IV U18467 ( .A(n18699), .Z(n18698) );
  XOR U18468 ( .A(n18700), .B(n18701), .Z(n18693) );
  ANDN U18469 ( .A(n18702), .B(n18564), .Z(n18701) );
  XNOR U18470 ( .A(n18700), .B(n18703), .Z(n18564) );
  XNOR U18471 ( .A(n18700), .B(n18562), .Z(n18702) );
  XOR U18472 ( .A(n18704), .B(n18705), .Z(n18562) );
  IV U18473 ( .A(n18706), .Z(n18705) );
  XOR U18474 ( .A(n18707), .B(n18708), .Z(n18700) );
  ANDN U18475 ( .A(n18709), .B(n18570), .Z(n18708) );
  XNOR U18476 ( .A(n18707), .B(n18710), .Z(n18570) );
  XNOR U18477 ( .A(n18707), .B(n18568), .Z(n18709) );
  XOR U18478 ( .A(n18711), .B(n18712), .Z(n18568) );
  IV U18479 ( .A(n18713), .Z(n18712) );
  XOR U18480 ( .A(n18714), .B(n18715), .Z(n18707) );
  NANDN U18481 ( .B(n18574), .A(n18716), .Z(n18714) );
  XOR U18482 ( .A(n18715), .B(n18572), .Z(n18716) );
  XOR U18483 ( .A(n18717), .B(n18718), .Z(n18572) );
  IV U18484 ( .A(n18719), .Z(n18718) );
  XNOR U18485 ( .A(n18720), .B(n18715), .Z(n18574) );
  OR U18486 ( .A(n12963), .B(n12964), .Z(n18715) );
  XOR U18487 ( .A(n18721), .B(n18722), .Z(n12963) );
  IV U18488 ( .A(n18723), .Z(n18722) );
  NAND U18489 ( .A(n16747), .B(n18675), .Z(n18720) );
  XOR U18490 ( .A(n16722), .B(n18724), .Z(n16716) );
  IV U18491 ( .A(n16721), .Z(n18724) );
  XNOR U18492 ( .A(n16718), .B(n16849), .Z(n16721) );
  AND U18493 ( .A(n18836), .B(n14041), .Z(n16849) );
  XOR U18494 ( .A(n18725), .B(n18726), .Z(n16718) );
  ANDN U18495 ( .A(n18727), .B(n18581), .Z(n18726) );
  XNOR U18496 ( .A(n18725), .B(n16893), .Z(n18581) );
  AND U18497 ( .A(n18836), .B(n14228), .Z(n16893) );
  XNOR U18498 ( .A(n18725), .B(n18579), .Z(n18727) );
  XOR U18499 ( .A(n18728), .B(n18729), .Z(n18579) );
  IV U18500 ( .A(n18730), .Z(n18729) );
  XOR U18501 ( .A(n18731), .B(n18732), .Z(n18725) );
  ANDN U18502 ( .A(n18733), .B(n18587), .Z(n18732) );
  XNOR U18503 ( .A(n18731), .B(n16947), .Z(n18587) );
  AND U18504 ( .A(n18836), .B(n14441), .Z(n16947) );
  XNOR U18505 ( .A(n18731), .B(n18585), .Z(n18733) );
  XOR U18506 ( .A(n18734), .B(n18735), .Z(n18585) );
  IV U18507 ( .A(n18736), .Z(n18735) );
  XOR U18508 ( .A(n18737), .B(n18738), .Z(n18731) );
  ANDN U18509 ( .A(n18739), .B(n18593), .Z(n18738) );
  XNOR U18510 ( .A(n18737), .B(n17008), .Z(n18593) );
  AND U18511 ( .A(n18836), .B(n14680), .Z(n17008) );
  XNOR U18512 ( .A(n18737), .B(n18591), .Z(n18739) );
  XOR U18513 ( .A(n18740), .B(n18741), .Z(n18591) );
  IV U18514 ( .A(n18742), .Z(n18741) );
  XOR U18515 ( .A(n18743), .B(n18744), .Z(n18737) );
  ANDN U18516 ( .A(n18745), .B(n18599), .Z(n18744) );
  XNOR U18517 ( .A(n18743), .B(n17076), .Z(n18599) );
  AND U18518 ( .A(n18836), .B(n14945), .Z(n17076) );
  XNOR U18519 ( .A(n18743), .B(n18597), .Z(n18745) );
  XOR U18520 ( .A(n18746), .B(n18747), .Z(n18597) );
  IV U18521 ( .A(n18748), .Z(n18747) );
  XOR U18522 ( .A(n18749), .B(n18750), .Z(n18743) );
  ANDN U18523 ( .A(n18751), .B(n18605), .Z(n18750) );
  XNOR U18524 ( .A(n18749), .B(n17151), .Z(n18605) );
  AND U18525 ( .A(n18836), .B(n15236), .Z(n17151) );
  XNOR U18526 ( .A(n18749), .B(n18603), .Z(n18751) );
  XOR U18527 ( .A(n18752), .B(n18753), .Z(n18603) );
  IV U18528 ( .A(n18754), .Z(n18753) );
  XOR U18529 ( .A(n18755), .B(n18756), .Z(n18749) );
  ANDN U18530 ( .A(n18757), .B(n18611), .Z(n18756) );
  XNOR U18531 ( .A(n18755), .B(n17233), .Z(n18611) );
  AND U18532 ( .A(n18836), .B(n15553), .Z(n17233) );
  XNOR U18533 ( .A(n18755), .B(n18609), .Z(n18757) );
  XOR U18534 ( .A(n18758), .B(n18759), .Z(n18609) );
  IV U18535 ( .A(n18760), .Z(n18759) );
  XOR U18536 ( .A(n18761), .B(n18762), .Z(n18755) );
  ANDN U18537 ( .A(n18763), .B(n18617), .Z(n18762) );
  XNOR U18538 ( .A(n18761), .B(n17322), .Z(n18617) );
  AND U18539 ( .A(n18836), .B(n15896), .Z(n17322) );
  XNOR U18540 ( .A(n18761), .B(n18615), .Z(n18763) );
  XOR U18541 ( .A(n18764), .B(n18765), .Z(n18615) );
  IV U18542 ( .A(n18766), .Z(n18765) );
  XOR U18543 ( .A(n18767), .B(n18768), .Z(n18761) );
  ANDN U18544 ( .A(n18769), .B(n18623), .Z(n18768) );
  XNOR U18545 ( .A(n18767), .B(n17418), .Z(n18623) );
  AND U18546 ( .A(n18836), .B(n16265), .Z(n17418) );
  XNOR U18547 ( .A(n18767), .B(n18621), .Z(n18769) );
  XOR U18548 ( .A(n18770), .B(n18771), .Z(n18621) );
  IV U18549 ( .A(n18772), .Z(n18771) );
  XOR U18550 ( .A(n18773), .B(n18774), .Z(n18767) );
  ANDN U18551 ( .A(n18775), .B(n18629), .Z(n18774) );
  XNOR U18552 ( .A(n18773), .B(n17521), .Z(n18629) );
  AND U18553 ( .A(n18836), .B(n16657), .Z(n17521) );
  XNOR U18554 ( .A(n18773), .B(n18627), .Z(n18775) );
  XOR U18555 ( .A(n18776), .B(n18777), .Z(n18627) );
  IV U18556 ( .A(n18778), .Z(n18777) );
  XOR U18557 ( .A(n18779), .B(n18780), .Z(n18773) );
  ANDN U18558 ( .A(n18781), .B(n18635), .Z(n18780) );
  XNOR U18559 ( .A(n18779), .B(n17630), .Z(n18635) );
  AND U18560 ( .A(n18836), .B(n17567), .Z(n17630) );
  XNOR U18561 ( .A(n18779), .B(n18633), .Z(n18781) );
  XOR U18562 ( .A(n18782), .B(n18783), .Z(n18633) );
  IV U18563 ( .A(n18784), .Z(n18783) );
  XOR U18564 ( .A(n18785), .B(n18786), .Z(n18779) );
  ANDN U18565 ( .A(n18787), .B(n18641), .Z(n18786) );
  XNOR U18566 ( .A(n18785), .B(n17744), .Z(n18641) );
  AND U18567 ( .A(n18836), .B(n17688), .Z(n17744) );
  XNOR U18568 ( .A(n18785), .B(n18639), .Z(n18787) );
  XOR U18569 ( .A(n18788), .B(n18789), .Z(n18639) );
  IV U18570 ( .A(n18790), .Z(n18789) );
  XOR U18571 ( .A(n18791), .B(n18792), .Z(n18785) );
  ANDN U18572 ( .A(n18793), .B(n18647), .Z(n18792) );
  XNOR U18573 ( .A(n18791), .B(n17863), .Z(n18647) );
  AND U18574 ( .A(n18836), .B(n17814), .Z(n17863) );
  XNOR U18575 ( .A(n18791), .B(n18645), .Z(n18793) );
  XOR U18576 ( .A(n18794), .B(n18795), .Z(n18645) );
  IV U18577 ( .A(n18796), .Z(n18795) );
  XOR U18578 ( .A(n18797), .B(n18798), .Z(n18791) );
  ANDN U18579 ( .A(n18799), .B(n18653), .Z(n18798) );
  XNOR U18580 ( .A(n18797), .B(n17987), .Z(n18653) );
  AND U18581 ( .A(n18836), .B(n17945), .Z(n17987) );
  XNOR U18582 ( .A(n18797), .B(n18651), .Z(n18799) );
  XOR U18583 ( .A(n18800), .B(n18801), .Z(n18651) );
  IV U18584 ( .A(n18802), .Z(n18801) );
  XOR U18585 ( .A(n18803), .B(n18804), .Z(n18797) );
  ANDN U18586 ( .A(n18805), .B(n18659), .Z(n18804) );
  XNOR U18587 ( .A(n18803), .B(n18116), .Z(n18659) );
  AND U18588 ( .A(n18836), .B(n18081), .Z(n18116) );
  XNOR U18589 ( .A(n18803), .B(n18657), .Z(n18805) );
  XOR U18590 ( .A(n18806), .B(n18807), .Z(n18657) );
  IV U18591 ( .A(n18808), .Z(n18807) );
  XOR U18592 ( .A(n18809), .B(n18810), .Z(n18803) );
  ANDN U18593 ( .A(n18811), .B(n18665), .Z(n18810) );
  XNOR U18594 ( .A(n18809), .B(n18250), .Z(n18665) );
  AND U18595 ( .A(n18836), .B(n18222), .Z(n18250) );
  XNOR U18596 ( .A(n18809), .B(n18663), .Z(n18811) );
  XOR U18597 ( .A(n18812), .B(n18813), .Z(n18663) );
  IV U18598 ( .A(n18814), .Z(n18813) );
  XOR U18599 ( .A(n18815), .B(n18816), .Z(n18809) );
  ANDN U18600 ( .A(n18817), .B(n18671), .Z(n18816) );
  XNOR U18601 ( .A(n18815), .B(n18389), .Z(n18671) );
  AND U18602 ( .A(n18836), .B(n18368), .Z(n18389) );
  XNOR U18603 ( .A(n18815), .B(n18669), .Z(n18817) );
  XOR U18604 ( .A(n18818), .B(n18819), .Z(n18669) );
  IV U18605 ( .A(n18820), .Z(n18819) );
  XOR U18606 ( .A(n18821), .B(n18822), .Z(n18815) );
  ANDN U18607 ( .A(n18823), .B(n18678), .Z(n18822) );
  XNOR U18608 ( .A(n18821), .B(n18533), .Z(n18678) );
  AND U18609 ( .A(n18836), .B(n18519), .Z(n18533) );
  XNOR U18610 ( .A(n18821), .B(n18676), .Z(n18823) );
  XOR U18611 ( .A(n18824), .B(n18825), .Z(n18676) );
  IV U18612 ( .A(n18826), .Z(n18825) );
  XOR U18613 ( .A(n18827), .B(n18828), .Z(n18821) );
  ANDN U18614 ( .A(n18829), .B(n18685), .Z(n18828) );
  XNOR U18615 ( .A(n18827), .B(n18682), .Z(n18685) );
  AND U18616 ( .A(n18836), .B(n18675), .Z(n18682) );
  XNOR U18617 ( .A(n18827), .B(n18683), .Z(n18829) );
  XOR U18618 ( .A(n18830), .B(n18831), .Z(n18683) );
  IV U18619 ( .A(n18832), .Z(n18831) );
  XOR U18620 ( .A(n18833), .B(n18834), .Z(n18827) );
  ANDN U18621 ( .A(n18835), .B(n18692), .Z(n18834) );
  XNOR U18622 ( .A(n18833), .B(n18836), .Z(n18692) );
  XNOR U18623 ( .A(n18833), .B(n18690), .Z(n18835) );
  XOR U18624 ( .A(n18837), .B(n18838), .Z(n18690) );
  IV U18625 ( .A(n18839), .Z(n18838) );
  XOR U18626 ( .A(n18840), .B(n18841), .Z(n18833) );
  ANDN U18627 ( .A(n18842), .B(n18699), .Z(n18841) );
  XNOR U18628 ( .A(n18840), .B(n18843), .Z(n18699) );
  XNOR U18629 ( .A(n18840), .B(n18697), .Z(n18842) );
  XOR U18630 ( .A(n18844), .B(n18845), .Z(n18697) );
  IV U18631 ( .A(n18846), .Z(n18845) );
  XOR U18632 ( .A(n18847), .B(n18848), .Z(n18840) );
  ANDN U18633 ( .A(n18849), .B(n18706), .Z(n18848) );
  XNOR U18634 ( .A(n18847), .B(n18850), .Z(n18706) );
  XNOR U18635 ( .A(n18847), .B(n18704), .Z(n18849) );
  XOR U18636 ( .A(n18851), .B(n18852), .Z(n18704) );
  IV U18637 ( .A(n18853), .Z(n18852) );
  XOR U18638 ( .A(n18854), .B(n18855), .Z(n18847) );
  ANDN U18639 ( .A(n18856), .B(n18713), .Z(n18855) );
  XNOR U18640 ( .A(n18854), .B(n18857), .Z(n18713) );
  XNOR U18641 ( .A(n18854), .B(n18711), .Z(n18856) );
  XOR U18642 ( .A(n18858), .B(n18859), .Z(n18711) );
  IV U18643 ( .A(n18860), .Z(n18859) );
  XOR U18644 ( .A(n18861), .B(n18862), .Z(n18854) );
  ANDN U18645 ( .A(n18863), .B(n18719), .Z(n18862) );
  XNOR U18646 ( .A(n18861), .B(n18864), .Z(n18719) );
  XNOR U18647 ( .A(n18861), .B(n18717), .Z(n18863) );
  XOR U18648 ( .A(n18865), .B(n18866), .Z(n18717) );
  IV U18649 ( .A(n18867), .Z(n18866) );
  XOR U18650 ( .A(n18868), .B(n18869), .Z(n18861) );
  NANDN U18651 ( .B(n18723), .A(n18870), .Z(n18868) );
  XOR U18652 ( .A(n18869), .B(n18721), .Z(n18870) );
  XOR U18653 ( .A(n18871), .B(n18872), .Z(n18721) );
  IV U18654 ( .A(n18873), .Z(n18872) );
  XNOR U18655 ( .A(n18874), .B(n18869), .Z(n18723) );
  OR U18656 ( .A(n13055), .B(n13056), .Z(n18869) );
  XOR U18657 ( .A(n18875), .B(n18876), .Z(n13055) );
  IV U18658 ( .A(n18877), .Z(n18876) );
  NAND U18659 ( .A(n16747), .B(n18836), .Z(n18874) );
  XOR U18660 ( .A(n16728), .B(n18878), .Z(n16722) );
  IV U18661 ( .A(n16727), .Z(n18878) );
  XNOR U18662 ( .A(n16724), .B(n16816), .Z(n16727) );
  AND U18663 ( .A(n19002), .B(n13880), .Z(n16816) );
  XOR U18664 ( .A(n18879), .B(n18880), .Z(n16724) );
  ANDN U18665 ( .A(n18881), .B(n18730), .Z(n18880) );
  XNOR U18666 ( .A(n18879), .B(n16853), .Z(n18730) );
  AND U18667 ( .A(n19002), .B(n14041), .Z(n16853) );
  XNOR U18668 ( .A(n18879), .B(n18728), .Z(n18881) );
  XOR U18669 ( .A(n18882), .B(n18883), .Z(n18728) );
  IV U18670 ( .A(n18884), .Z(n18883) );
  XOR U18671 ( .A(n18885), .B(n18886), .Z(n18879) );
  ANDN U18672 ( .A(n18887), .B(n18736), .Z(n18886) );
  XNOR U18673 ( .A(n18885), .B(n16900), .Z(n18736) );
  AND U18674 ( .A(n19002), .B(n14228), .Z(n16900) );
  XNOR U18675 ( .A(n18885), .B(n18734), .Z(n18887) );
  XOR U18676 ( .A(n18888), .B(n18889), .Z(n18734) );
  IV U18677 ( .A(n18890), .Z(n18889) );
  XOR U18678 ( .A(n18891), .B(n18892), .Z(n18885) );
  ANDN U18679 ( .A(n18893), .B(n18742), .Z(n18892) );
  XNOR U18680 ( .A(n18891), .B(n16954), .Z(n18742) );
  AND U18681 ( .A(n19002), .B(n14441), .Z(n16954) );
  XNOR U18682 ( .A(n18891), .B(n18740), .Z(n18893) );
  XOR U18683 ( .A(n18894), .B(n18895), .Z(n18740) );
  IV U18684 ( .A(n18896), .Z(n18895) );
  XOR U18685 ( .A(n18897), .B(n18898), .Z(n18891) );
  ANDN U18686 ( .A(n18899), .B(n18748), .Z(n18898) );
  XNOR U18687 ( .A(n18897), .B(n17015), .Z(n18748) );
  AND U18688 ( .A(n19002), .B(n14680), .Z(n17015) );
  XNOR U18689 ( .A(n18897), .B(n18746), .Z(n18899) );
  XOR U18690 ( .A(n18900), .B(n18901), .Z(n18746) );
  IV U18691 ( .A(n18902), .Z(n18901) );
  XOR U18692 ( .A(n18903), .B(n18904), .Z(n18897) );
  ANDN U18693 ( .A(n18905), .B(n18754), .Z(n18904) );
  XNOR U18694 ( .A(n18903), .B(n17083), .Z(n18754) );
  AND U18695 ( .A(n19002), .B(n14945), .Z(n17083) );
  XNOR U18696 ( .A(n18903), .B(n18752), .Z(n18905) );
  XOR U18697 ( .A(n18906), .B(n18907), .Z(n18752) );
  IV U18698 ( .A(n18908), .Z(n18907) );
  XOR U18699 ( .A(n18909), .B(n18910), .Z(n18903) );
  ANDN U18700 ( .A(n18911), .B(n18760), .Z(n18910) );
  XNOR U18701 ( .A(n18909), .B(n17158), .Z(n18760) );
  AND U18702 ( .A(n19002), .B(n15236), .Z(n17158) );
  XNOR U18703 ( .A(n18909), .B(n18758), .Z(n18911) );
  XOR U18704 ( .A(n18912), .B(n18913), .Z(n18758) );
  IV U18705 ( .A(n18914), .Z(n18913) );
  XOR U18706 ( .A(n18915), .B(n18916), .Z(n18909) );
  ANDN U18707 ( .A(n18917), .B(n18766), .Z(n18916) );
  XNOR U18708 ( .A(n18915), .B(n17240), .Z(n18766) );
  AND U18709 ( .A(n19002), .B(n15553), .Z(n17240) );
  XNOR U18710 ( .A(n18915), .B(n18764), .Z(n18917) );
  XOR U18711 ( .A(n18918), .B(n18919), .Z(n18764) );
  IV U18712 ( .A(n18920), .Z(n18919) );
  XOR U18713 ( .A(n18921), .B(n18922), .Z(n18915) );
  ANDN U18714 ( .A(n18923), .B(n18772), .Z(n18922) );
  XNOR U18715 ( .A(n18921), .B(n17329), .Z(n18772) );
  AND U18716 ( .A(n19002), .B(n15896), .Z(n17329) );
  XNOR U18717 ( .A(n18921), .B(n18770), .Z(n18923) );
  XOR U18718 ( .A(n18924), .B(n18925), .Z(n18770) );
  IV U18719 ( .A(n18926), .Z(n18925) );
  XOR U18720 ( .A(n18927), .B(n18928), .Z(n18921) );
  ANDN U18721 ( .A(n18929), .B(n18778), .Z(n18928) );
  XNOR U18722 ( .A(n18927), .B(n17425), .Z(n18778) );
  AND U18723 ( .A(n19002), .B(n16265), .Z(n17425) );
  XNOR U18724 ( .A(n18927), .B(n18776), .Z(n18929) );
  XOR U18725 ( .A(n18930), .B(n18931), .Z(n18776) );
  IV U18726 ( .A(n18932), .Z(n18931) );
  XOR U18727 ( .A(n18933), .B(n18934), .Z(n18927) );
  ANDN U18728 ( .A(n18935), .B(n18784), .Z(n18934) );
  XNOR U18729 ( .A(n18933), .B(n17528), .Z(n18784) );
  AND U18730 ( .A(n19002), .B(n16657), .Z(n17528) );
  XNOR U18731 ( .A(n18933), .B(n18782), .Z(n18935) );
  XOR U18732 ( .A(n18936), .B(n18937), .Z(n18782) );
  IV U18733 ( .A(n18938), .Z(n18937) );
  XOR U18734 ( .A(n18939), .B(n18940), .Z(n18933) );
  ANDN U18735 ( .A(n18941), .B(n18790), .Z(n18940) );
  XNOR U18736 ( .A(n18939), .B(n17637), .Z(n18790) );
  AND U18737 ( .A(n19002), .B(n17567), .Z(n17637) );
  XNOR U18738 ( .A(n18939), .B(n18788), .Z(n18941) );
  XOR U18739 ( .A(n18942), .B(n18943), .Z(n18788) );
  IV U18740 ( .A(n18944), .Z(n18943) );
  XOR U18741 ( .A(n18945), .B(n18946), .Z(n18939) );
  ANDN U18742 ( .A(n18947), .B(n18796), .Z(n18946) );
  XNOR U18743 ( .A(n18945), .B(n17751), .Z(n18796) );
  AND U18744 ( .A(n19002), .B(n17688), .Z(n17751) );
  XNOR U18745 ( .A(n18945), .B(n18794), .Z(n18947) );
  XOR U18746 ( .A(n18948), .B(n18949), .Z(n18794) );
  IV U18747 ( .A(n18950), .Z(n18949) );
  XOR U18748 ( .A(n18951), .B(n18952), .Z(n18945) );
  ANDN U18749 ( .A(n18953), .B(n18802), .Z(n18952) );
  XNOR U18750 ( .A(n18951), .B(n17870), .Z(n18802) );
  AND U18751 ( .A(n19002), .B(n17814), .Z(n17870) );
  XNOR U18752 ( .A(n18951), .B(n18800), .Z(n18953) );
  XOR U18753 ( .A(n18954), .B(n18955), .Z(n18800) );
  IV U18754 ( .A(n18956), .Z(n18955) );
  XOR U18755 ( .A(n18957), .B(n18958), .Z(n18951) );
  ANDN U18756 ( .A(n18959), .B(n18808), .Z(n18958) );
  XNOR U18757 ( .A(n18957), .B(n17994), .Z(n18808) );
  AND U18758 ( .A(n19002), .B(n17945), .Z(n17994) );
  XNOR U18759 ( .A(n18957), .B(n18806), .Z(n18959) );
  XOR U18760 ( .A(n18960), .B(n18961), .Z(n18806) );
  IV U18761 ( .A(n18962), .Z(n18961) );
  XOR U18762 ( .A(n18963), .B(n18964), .Z(n18957) );
  ANDN U18763 ( .A(n18965), .B(n18814), .Z(n18964) );
  XNOR U18764 ( .A(n18963), .B(n18123), .Z(n18814) );
  AND U18765 ( .A(n19002), .B(n18081), .Z(n18123) );
  XNOR U18766 ( .A(n18963), .B(n18812), .Z(n18965) );
  XOR U18767 ( .A(n18966), .B(n18967), .Z(n18812) );
  IV U18768 ( .A(n18968), .Z(n18967) );
  XOR U18769 ( .A(n18969), .B(n18970), .Z(n18963) );
  ANDN U18770 ( .A(n18971), .B(n18820), .Z(n18970) );
  XNOR U18771 ( .A(n18969), .B(n18257), .Z(n18820) );
  AND U18772 ( .A(n19002), .B(n18222), .Z(n18257) );
  XNOR U18773 ( .A(n18969), .B(n18818), .Z(n18971) );
  XOR U18774 ( .A(n18972), .B(n18973), .Z(n18818) );
  IV U18775 ( .A(n18974), .Z(n18973) );
  XOR U18776 ( .A(n18975), .B(n18976), .Z(n18969) );
  ANDN U18777 ( .A(n18977), .B(n18826), .Z(n18976) );
  XNOR U18778 ( .A(n18975), .B(n18396), .Z(n18826) );
  AND U18779 ( .A(n19002), .B(n18368), .Z(n18396) );
  XNOR U18780 ( .A(n18975), .B(n18824), .Z(n18977) );
  XOR U18781 ( .A(n18978), .B(n18979), .Z(n18824) );
  IV U18782 ( .A(n18980), .Z(n18979) );
  XOR U18783 ( .A(n18981), .B(n18982), .Z(n18975) );
  ANDN U18784 ( .A(n18983), .B(n18832), .Z(n18982) );
  XNOR U18785 ( .A(n18981), .B(n18540), .Z(n18832) );
  AND U18786 ( .A(n19002), .B(n18519), .Z(n18540) );
  XNOR U18787 ( .A(n18981), .B(n18830), .Z(n18983) );
  XOR U18788 ( .A(n18984), .B(n18985), .Z(n18830) );
  IV U18789 ( .A(n18986), .Z(n18985) );
  XOR U18790 ( .A(n18987), .B(n18988), .Z(n18981) );
  ANDN U18791 ( .A(n18989), .B(n18839), .Z(n18988) );
  XNOR U18792 ( .A(n18987), .B(n18689), .Z(n18839) );
  AND U18793 ( .A(n19002), .B(n18675), .Z(n18689) );
  XNOR U18794 ( .A(n18987), .B(n18837), .Z(n18989) );
  XOR U18795 ( .A(n18990), .B(n18991), .Z(n18837) );
  IV U18796 ( .A(n18992), .Z(n18991) );
  XOR U18797 ( .A(n18993), .B(n18994), .Z(n18987) );
  ANDN U18798 ( .A(n18995), .B(n18846), .Z(n18994) );
  XNOR U18799 ( .A(n18993), .B(n18843), .Z(n18846) );
  AND U18800 ( .A(n19002), .B(n18836), .Z(n18843) );
  XNOR U18801 ( .A(n18993), .B(n18844), .Z(n18995) );
  XOR U18802 ( .A(n18996), .B(n18997), .Z(n18844) );
  IV U18803 ( .A(n18998), .Z(n18997) );
  XOR U18804 ( .A(n18999), .B(n19000), .Z(n18993) );
  ANDN U18805 ( .A(n19001), .B(n18853), .Z(n19000) );
  XNOR U18806 ( .A(n18999), .B(n19002), .Z(n18853) );
  XNOR U18807 ( .A(n18999), .B(n18851), .Z(n19001) );
  XOR U18808 ( .A(n19003), .B(n19004), .Z(n18851) );
  IV U18809 ( .A(n19005), .Z(n19004) );
  XOR U18810 ( .A(n19006), .B(n19007), .Z(n18999) );
  ANDN U18811 ( .A(n19008), .B(n18860), .Z(n19007) );
  XNOR U18812 ( .A(n19006), .B(n19009), .Z(n18860) );
  XNOR U18813 ( .A(n19006), .B(n18858), .Z(n19008) );
  XOR U18814 ( .A(n19010), .B(n19011), .Z(n18858) );
  IV U18815 ( .A(n19012), .Z(n19011) );
  XOR U18816 ( .A(n19013), .B(n19014), .Z(n19006) );
  ANDN U18817 ( .A(n19015), .B(n18867), .Z(n19014) );
  XNOR U18818 ( .A(n19013), .B(n19016), .Z(n18867) );
  XNOR U18819 ( .A(n19013), .B(n18865), .Z(n19015) );
  XOR U18820 ( .A(n19017), .B(n19018), .Z(n18865) );
  IV U18821 ( .A(n19019), .Z(n19018) );
  XOR U18822 ( .A(n19020), .B(n19021), .Z(n19013) );
  ANDN U18823 ( .A(n19022), .B(n18873), .Z(n19021) );
  XNOR U18824 ( .A(n19020), .B(n19023), .Z(n18873) );
  XNOR U18825 ( .A(n19020), .B(n18871), .Z(n19022) );
  XOR U18826 ( .A(n19024), .B(n19025), .Z(n18871) );
  IV U18827 ( .A(n19026), .Z(n19025) );
  XOR U18828 ( .A(n19027), .B(n19028), .Z(n19020) );
  NANDN U18829 ( .B(n18877), .A(n19029), .Z(n19027) );
  XOR U18830 ( .A(n19028), .B(n18875), .Z(n19029) );
  XOR U18831 ( .A(n19030), .B(n19031), .Z(n18875) );
  IV U18832 ( .A(n19032), .Z(n19031) );
  XNOR U18833 ( .A(n19033), .B(n19028), .Z(n18877) );
  OR U18834 ( .A(n13134), .B(n13135), .Z(n19028) );
  XOR U18835 ( .A(n19034), .B(n19035), .Z(n13134) );
  IV U18836 ( .A(n19036), .Z(n19035) );
  NAND U18837 ( .A(n16747), .B(n19002), .Z(n19033) );
  XOR U18838 ( .A(n16734), .B(n19037), .Z(n16728) );
  IV U18839 ( .A(n16733), .Z(n19037) );
  XNOR U18840 ( .A(n16730), .B(n16790), .Z(n16733) );
  AND U18841 ( .A(n19173), .B(n13745), .Z(n16790) );
  XOR U18842 ( .A(n19038), .B(n19039), .Z(n16730) );
  ANDN U18843 ( .A(n19040), .B(n18884), .Z(n19039) );
  XNOR U18844 ( .A(n19038), .B(n16820), .Z(n18884) );
  AND U18845 ( .A(n19173), .B(n13880), .Z(n16820) );
  XNOR U18846 ( .A(n19038), .B(n18882), .Z(n19040) );
  XOR U18847 ( .A(n19041), .B(n19042), .Z(n18882) );
  IV U18848 ( .A(n19043), .Z(n19042) );
  XOR U18849 ( .A(n19044), .B(n19045), .Z(n19038) );
  ANDN U18850 ( .A(n19046), .B(n18890), .Z(n19045) );
  XNOR U18851 ( .A(n19044), .B(n16860), .Z(n18890) );
  AND U18852 ( .A(n19173), .B(n14041), .Z(n16860) );
  XNOR U18853 ( .A(n19044), .B(n18888), .Z(n19046) );
  XOR U18854 ( .A(n19047), .B(n19048), .Z(n18888) );
  IV U18855 ( .A(n19049), .Z(n19048) );
  XOR U18856 ( .A(n19050), .B(n19051), .Z(n19044) );
  ANDN U18857 ( .A(n19052), .B(n18896), .Z(n19051) );
  XNOR U18858 ( .A(n19050), .B(n16907), .Z(n18896) );
  AND U18859 ( .A(n19173), .B(n14228), .Z(n16907) );
  XNOR U18860 ( .A(n19050), .B(n18894), .Z(n19052) );
  XOR U18861 ( .A(n19053), .B(n19054), .Z(n18894) );
  IV U18862 ( .A(n19055), .Z(n19054) );
  XOR U18863 ( .A(n19056), .B(n19057), .Z(n19050) );
  ANDN U18864 ( .A(n19058), .B(n18902), .Z(n19057) );
  XNOR U18865 ( .A(n19056), .B(n16961), .Z(n18902) );
  AND U18866 ( .A(n19173), .B(n14441), .Z(n16961) );
  XNOR U18867 ( .A(n19056), .B(n18900), .Z(n19058) );
  XOR U18868 ( .A(n19059), .B(n19060), .Z(n18900) );
  IV U18869 ( .A(n19061), .Z(n19060) );
  XOR U18870 ( .A(n19062), .B(n19063), .Z(n19056) );
  ANDN U18871 ( .A(n19064), .B(n18908), .Z(n19063) );
  XNOR U18872 ( .A(n19062), .B(n17022), .Z(n18908) );
  AND U18873 ( .A(n19173), .B(n14680), .Z(n17022) );
  XNOR U18874 ( .A(n19062), .B(n18906), .Z(n19064) );
  XOR U18875 ( .A(n19065), .B(n19066), .Z(n18906) );
  IV U18876 ( .A(n19067), .Z(n19066) );
  XOR U18877 ( .A(n19068), .B(n19069), .Z(n19062) );
  ANDN U18878 ( .A(n19070), .B(n18914), .Z(n19069) );
  XNOR U18879 ( .A(n19068), .B(n17090), .Z(n18914) );
  AND U18880 ( .A(n19173), .B(n14945), .Z(n17090) );
  XNOR U18881 ( .A(n19068), .B(n18912), .Z(n19070) );
  XOR U18882 ( .A(n19071), .B(n19072), .Z(n18912) );
  IV U18883 ( .A(n19073), .Z(n19072) );
  XOR U18884 ( .A(n19074), .B(n19075), .Z(n19068) );
  ANDN U18885 ( .A(n19076), .B(n18920), .Z(n19075) );
  XNOR U18886 ( .A(n19074), .B(n17165), .Z(n18920) );
  AND U18887 ( .A(n19173), .B(n15236), .Z(n17165) );
  XNOR U18888 ( .A(n19074), .B(n18918), .Z(n19076) );
  XOR U18889 ( .A(n19077), .B(n19078), .Z(n18918) );
  IV U18890 ( .A(n19079), .Z(n19078) );
  XOR U18891 ( .A(n19080), .B(n19081), .Z(n19074) );
  ANDN U18892 ( .A(n19082), .B(n18926), .Z(n19081) );
  XNOR U18893 ( .A(n19080), .B(n17247), .Z(n18926) );
  AND U18894 ( .A(n19173), .B(n15553), .Z(n17247) );
  XNOR U18895 ( .A(n19080), .B(n18924), .Z(n19082) );
  XOR U18896 ( .A(n19083), .B(n19084), .Z(n18924) );
  IV U18897 ( .A(n19085), .Z(n19084) );
  XOR U18898 ( .A(n19086), .B(n19087), .Z(n19080) );
  ANDN U18899 ( .A(n19088), .B(n18932), .Z(n19087) );
  XNOR U18900 ( .A(n19086), .B(n17336), .Z(n18932) );
  AND U18901 ( .A(n19173), .B(n15896), .Z(n17336) );
  XNOR U18902 ( .A(n19086), .B(n18930), .Z(n19088) );
  XOR U18903 ( .A(n19089), .B(n19090), .Z(n18930) );
  IV U18904 ( .A(n19091), .Z(n19090) );
  XOR U18905 ( .A(n19092), .B(n19093), .Z(n19086) );
  ANDN U18906 ( .A(n19094), .B(n18938), .Z(n19093) );
  XNOR U18907 ( .A(n19092), .B(n17432), .Z(n18938) );
  AND U18908 ( .A(n19173), .B(n16265), .Z(n17432) );
  XNOR U18909 ( .A(n19092), .B(n18936), .Z(n19094) );
  XOR U18910 ( .A(n19095), .B(n19096), .Z(n18936) );
  IV U18911 ( .A(n19097), .Z(n19096) );
  XOR U18912 ( .A(n19098), .B(n19099), .Z(n19092) );
  ANDN U18913 ( .A(n19100), .B(n18944), .Z(n19099) );
  XNOR U18914 ( .A(n19098), .B(n17535), .Z(n18944) );
  AND U18915 ( .A(n19173), .B(n16657), .Z(n17535) );
  XNOR U18916 ( .A(n19098), .B(n18942), .Z(n19100) );
  XOR U18917 ( .A(n19101), .B(n19102), .Z(n18942) );
  IV U18918 ( .A(n19103), .Z(n19102) );
  XOR U18919 ( .A(n19104), .B(n19105), .Z(n19098) );
  ANDN U18920 ( .A(n19106), .B(n18950), .Z(n19105) );
  XNOR U18921 ( .A(n19104), .B(n17644), .Z(n18950) );
  AND U18922 ( .A(n19173), .B(n17567), .Z(n17644) );
  XNOR U18923 ( .A(n19104), .B(n18948), .Z(n19106) );
  XOR U18924 ( .A(n19107), .B(n19108), .Z(n18948) );
  IV U18925 ( .A(n19109), .Z(n19108) );
  XOR U18926 ( .A(n19110), .B(n19111), .Z(n19104) );
  ANDN U18927 ( .A(n19112), .B(n18956), .Z(n19111) );
  XNOR U18928 ( .A(n19110), .B(n17758), .Z(n18956) );
  AND U18929 ( .A(n19173), .B(n17688), .Z(n17758) );
  XNOR U18930 ( .A(n19110), .B(n18954), .Z(n19112) );
  XOR U18931 ( .A(n19113), .B(n19114), .Z(n18954) );
  IV U18932 ( .A(n19115), .Z(n19114) );
  XOR U18933 ( .A(n19116), .B(n19117), .Z(n19110) );
  ANDN U18934 ( .A(n19118), .B(n18962), .Z(n19117) );
  XNOR U18935 ( .A(n19116), .B(n17877), .Z(n18962) );
  AND U18936 ( .A(n19173), .B(n17814), .Z(n17877) );
  XNOR U18937 ( .A(n19116), .B(n18960), .Z(n19118) );
  XOR U18938 ( .A(n19119), .B(n19120), .Z(n18960) );
  IV U18939 ( .A(n19121), .Z(n19120) );
  XOR U18940 ( .A(n19122), .B(n19123), .Z(n19116) );
  ANDN U18941 ( .A(n19124), .B(n18968), .Z(n19123) );
  XNOR U18942 ( .A(n19122), .B(n18001), .Z(n18968) );
  AND U18943 ( .A(n19173), .B(n17945), .Z(n18001) );
  XNOR U18944 ( .A(n19122), .B(n18966), .Z(n19124) );
  XOR U18945 ( .A(n19125), .B(n19126), .Z(n18966) );
  IV U18946 ( .A(n19127), .Z(n19126) );
  XOR U18947 ( .A(n19128), .B(n19129), .Z(n19122) );
  ANDN U18948 ( .A(n19130), .B(n18974), .Z(n19129) );
  XNOR U18949 ( .A(n19128), .B(n18130), .Z(n18974) );
  AND U18950 ( .A(n19173), .B(n18081), .Z(n18130) );
  XNOR U18951 ( .A(n19128), .B(n18972), .Z(n19130) );
  XOR U18952 ( .A(n19131), .B(n19132), .Z(n18972) );
  IV U18953 ( .A(n19133), .Z(n19132) );
  XOR U18954 ( .A(n19134), .B(n19135), .Z(n19128) );
  ANDN U18955 ( .A(n19136), .B(n18980), .Z(n19135) );
  XNOR U18956 ( .A(n19134), .B(n18264), .Z(n18980) );
  AND U18957 ( .A(n19173), .B(n18222), .Z(n18264) );
  XNOR U18958 ( .A(n19134), .B(n18978), .Z(n19136) );
  XOR U18959 ( .A(n19137), .B(n19138), .Z(n18978) );
  IV U18960 ( .A(n19139), .Z(n19138) );
  XOR U18961 ( .A(n19140), .B(n19141), .Z(n19134) );
  ANDN U18962 ( .A(n19142), .B(n18986), .Z(n19141) );
  XNOR U18963 ( .A(n19140), .B(n18403), .Z(n18986) );
  AND U18964 ( .A(n19173), .B(n18368), .Z(n18403) );
  XNOR U18965 ( .A(n19140), .B(n18984), .Z(n19142) );
  XOR U18966 ( .A(n19143), .B(n19144), .Z(n18984) );
  IV U18967 ( .A(n19145), .Z(n19144) );
  XOR U18968 ( .A(n19146), .B(n19147), .Z(n19140) );
  ANDN U18969 ( .A(n19148), .B(n18992), .Z(n19147) );
  XNOR U18970 ( .A(n19146), .B(n18547), .Z(n18992) );
  AND U18971 ( .A(n19173), .B(n18519), .Z(n18547) );
  XNOR U18972 ( .A(n19146), .B(n18990), .Z(n19148) );
  XOR U18973 ( .A(n19149), .B(n19150), .Z(n18990) );
  IV U18974 ( .A(n19151), .Z(n19150) );
  XOR U18975 ( .A(n19152), .B(n19153), .Z(n19146) );
  ANDN U18976 ( .A(n19154), .B(n18998), .Z(n19153) );
  XNOR U18977 ( .A(n19152), .B(n18696), .Z(n18998) );
  AND U18978 ( .A(n19173), .B(n18675), .Z(n18696) );
  XNOR U18979 ( .A(n19152), .B(n18996), .Z(n19154) );
  XOR U18980 ( .A(n19155), .B(n19156), .Z(n18996) );
  IV U18981 ( .A(n19157), .Z(n19156) );
  XOR U18982 ( .A(n19158), .B(n19159), .Z(n19152) );
  ANDN U18983 ( .A(n19160), .B(n19005), .Z(n19159) );
  XNOR U18984 ( .A(n19158), .B(n18850), .Z(n19005) );
  AND U18985 ( .A(n19173), .B(n18836), .Z(n18850) );
  XNOR U18986 ( .A(n19158), .B(n19003), .Z(n19160) );
  XOR U18987 ( .A(n19161), .B(n19162), .Z(n19003) );
  IV U18988 ( .A(n19163), .Z(n19162) );
  XOR U18989 ( .A(n19164), .B(n19165), .Z(n19158) );
  ANDN U18990 ( .A(n19166), .B(n19012), .Z(n19165) );
  XNOR U18991 ( .A(n19164), .B(n19009), .Z(n19012) );
  AND U18992 ( .A(n19173), .B(n19002), .Z(n19009) );
  XNOR U18993 ( .A(n19164), .B(n19010), .Z(n19166) );
  XOR U18994 ( .A(n19167), .B(n19168), .Z(n19010) );
  IV U18995 ( .A(n19169), .Z(n19168) );
  XOR U18996 ( .A(n19170), .B(n19171), .Z(n19164) );
  ANDN U18997 ( .A(n19172), .B(n19019), .Z(n19171) );
  XNOR U18998 ( .A(n19170), .B(n19173), .Z(n19019) );
  XNOR U18999 ( .A(n19170), .B(n19017), .Z(n19172) );
  XOR U19000 ( .A(n19174), .B(n19175), .Z(n19017) );
  IV U19001 ( .A(n19176), .Z(n19175) );
  XOR U19002 ( .A(n19177), .B(n19178), .Z(n19170) );
  ANDN U19003 ( .A(n19179), .B(n19026), .Z(n19178) );
  XNOR U19004 ( .A(n19177), .B(n19180), .Z(n19026) );
  XNOR U19005 ( .A(n19177), .B(n19024), .Z(n19179) );
  XOR U19006 ( .A(n19181), .B(n19182), .Z(n19024) );
  IV U19007 ( .A(n19183), .Z(n19182) );
  XOR U19008 ( .A(n19184), .B(n19185), .Z(n19177) );
  ANDN U19009 ( .A(n19186), .B(n19032), .Z(n19185) );
  XNOR U19010 ( .A(n19184), .B(n19187), .Z(n19032) );
  XNOR U19011 ( .A(n19184), .B(n19030), .Z(n19186) );
  XOR U19012 ( .A(n19188), .B(n19189), .Z(n19030) );
  IV U19013 ( .A(n19190), .Z(n19189) );
  XOR U19014 ( .A(n19191), .B(n19192), .Z(n19184) );
  NANDN U19015 ( .B(n19036), .A(n19193), .Z(n19191) );
  XOR U19016 ( .A(n19192), .B(n19034), .Z(n19193) );
  XOR U19017 ( .A(n19194), .B(n19195), .Z(n19034) );
  IV U19018 ( .A(n19196), .Z(n19195) );
  XNOR U19019 ( .A(n19197), .B(n19192), .Z(n19036) );
  OR U19020 ( .A(n13199), .B(n13200), .Z(n19192) );
  XOR U19021 ( .A(n19198), .B(n19199), .Z(n13199) );
  IV U19022 ( .A(n19200), .Z(n19199) );
  NAND U19023 ( .A(n16747), .B(n19173), .Z(n19197) );
  XOR U19024 ( .A(n16740), .B(n19201), .Z(n16734) );
  IV U19025 ( .A(n16739), .Z(n19201) );
  XNOR U19026 ( .A(n16736), .B(n16771), .Z(n16739) );
  AND U19027 ( .A(n19349), .B(n13636), .Z(n16771) );
  XOR U19028 ( .A(n19202), .B(n19203), .Z(n16736) );
  ANDN U19029 ( .A(n19204), .B(n19043), .Z(n19203) );
  XNOR U19030 ( .A(n19202), .B(n16794), .Z(n19043) );
  AND U19031 ( .A(n19349), .B(n13745), .Z(n16794) );
  XNOR U19032 ( .A(n19202), .B(n19041), .Z(n19204) );
  XOR U19033 ( .A(n19205), .B(n19206), .Z(n19041) );
  IV U19034 ( .A(n19207), .Z(n19206) );
  XOR U19035 ( .A(n19208), .B(n19209), .Z(n19202) );
  ANDN U19036 ( .A(n19210), .B(n19049), .Z(n19209) );
  XNOR U19037 ( .A(n19208), .B(n16827), .Z(n19049) );
  AND U19038 ( .A(n19349), .B(n13880), .Z(n16827) );
  XNOR U19039 ( .A(n19208), .B(n19047), .Z(n19210) );
  XOR U19040 ( .A(n19211), .B(n19212), .Z(n19047) );
  IV U19041 ( .A(n19213), .Z(n19212) );
  XOR U19042 ( .A(n19214), .B(n19215), .Z(n19208) );
  ANDN U19043 ( .A(n19216), .B(n19055), .Z(n19215) );
  XNOR U19044 ( .A(n19214), .B(n16867), .Z(n19055) );
  AND U19045 ( .A(n19349), .B(n14041), .Z(n16867) );
  XNOR U19046 ( .A(n19214), .B(n19053), .Z(n19216) );
  XOR U19047 ( .A(n19217), .B(n19218), .Z(n19053) );
  IV U19048 ( .A(n19219), .Z(n19218) );
  XOR U19049 ( .A(n19220), .B(n19221), .Z(n19214) );
  ANDN U19050 ( .A(n19222), .B(n19061), .Z(n19221) );
  XNOR U19051 ( .A(n19220), .B(n16914), .Z(n19061) );
  AND U19052 ( .A(n19349), .B(n14228), .Z(n16914) );
  XNOR U19053 ( .A(n19220), .B(n19059), .Z(n19222) );
  XOR U19054 ( .A(n19223), .B(n19224), .Z(n19059) );
  IV U19055 ( .A(n19225), .Z(n19224) );
  XOR U19056 ( .A(n19226), .B(n19227), .Z(n19220) );
  ANDN U19057 ( .A(n19228), .B(n19067), .Z(n19227) );
  XNOR U19058 ( .A(n19226), .B(n16968), .Z(n19067) );
  AND U19059 ( .A(n19349), .B(n14441), .Z(n16968) );
  XNOR U19060 ( .A(n19226), .B(n19065), .Z(n19228) );
  XOR U19061 ( .A(n19229), .B(n19230), .Z(n19065) );
  IV U19062 ( .A(n19231), .Z(n19230) );
  XOR U19063 ( .A(n19232), .B(n19233), .Z(n19226) );
  ANDN U19064 ( .A(n19234), .B(n19073), .Z(n19233) );
  XNOR U19065 ( .A(n19232), .B(n17029), .Z(n19073) );
  AND U19066 ( .A(n19349), .B(n14680), .Z(n17029) );
  XNOR U19067 ( .A(n19232), .B(n19071), .Z(n19234) );
  XOR U19068 ( .A(n19235), .B(n19236), .Z(n19071) );
  IV U19069 ( .A(n19237), .Z(n19236) );
  XOR U19070 ( .A(n19238), .B(n19239), .Z(n19232) );
  ANDN U19071 ( .A(n19240), .B(n19079), .Z(n19239) );
  XNOR U19072 ( .A(n19238), .B(n17097), .Z(n19079) );
  AND U19073 ( .A(n19349), .B(n14945), .Z(n17097) );
  XNOR U19074 ( .A(n19238), .B(n19077), .Z(n19240) );
  XOR U19075 ( .A(n19241), .B(n19242), .Z(n19077) );
  IV U19076 ( .A(n19243), .Z(n19242) );
  XOR U19077 ( .A(n19244), .B(n19245), .Z(n19238) );
  ANDN U19078 ( .A(n19246), .B(n19085), .Z(n19245) );
  XNOR U19079 ( .A(n19244), .B(n17172), .Z(n19085) );
  AND U19080 ( .A(n19349), .B(n15236), .Z(n17172) );
  XNOR U19081 ( .A(n19244), .B(n19083), .Z(n19246) );
  XOR U19082 ( .A(n19247), .B(n19248), .Z(n19083) );
  IV U19083 ( .A(n19249), .Z(n19248) );
  XOR U19084 ( .A(n19250), .B(n19251), .Z(n19244) );
  ANDN U19085 ( .A(n19252), .B(n19091), .Z(n19251) );
  XNOR U19086 ( .A(n19250), .B(n17254), .Z(n19091) );
  AND U19087 ( .A(n19349), .B(n15553), .Z(n17254) );
  XNOR U19088 ( .A(n19250), .B(n19089), .Z(n19252) );
  XOR U19089 ( .A(n19253), .B(n19254), .Z(n19089) );
  IV U19090 ( .A(n19255), .Z(n19254) );
  XOR U19091 ( .A(n19256), .B(n19257), .Z(n19250) );
  ANDN U19092 ( .A(n19258), .B(n19097), .Z(n19257) );
  XNOR U19093 ( .A(n19256), .B(n17343), .Z(n19097) );
  AND U19094 ( .A(n19349), .B(n15896), .Z(n17343) );
  XNOR U19095 ( .A(n19256), .B(n19095), .Z(n19258) );
  XOR U19096 ( .A(n19259), .B(n19260), .Z(n19095) );
  IV U19097 ( .A(n19261), .Z(n19260) );
  XOR U19098 ( .A(n19262), .B(n19263), .Z(n19256) );
  ANDN U19099 ( .A(n19264), .B(n19103), .Z(n19263) );
  XNOR U19100 ( .A(n19262), .B(n17439), .Z(n19103) );
  AND U19101 ( .A(n19349), .B(n16265), .Z(n17439) );
  XNOR U19102 ( .A(n19262), .B(n19101), .Z(n19264) );
  XOR U19103 ( .A(n19265), .B(n19266), .Z(n19101) );
  IV U19104 ( .A(n19267), .Z(n19266) );
  XOR U19105 ( .A(n19268), .B(n19269), .Z(n19262) );
  ANDN U19106 ( .A(n19270), .B(n19109), .Z(n19269) );
  XNOR U19107 ( .A(n19268), .B(n17542), .Z(n19109) );
  AND U19108 ( .A(n19349), .B(n16657), .Z(n17542) );
  XNOR U19109 ( .A(n19268), .B(n19107), .Z(n19270) );
  XOR U19110 ( .A(n19271), .B(n19272), .Z(n19107) );
  IV U19111 ( .A(n19273), .Z(n19272) );
  XOR U19112 ( .A(n19274), .B(n19275), .Z(n19268) );
  ANDN U19113 ( .A(n19276), .B(n19115), .Z(n19275) );
  XNOR U19114 ( .A(n19274), .B(n17651), .Z(n19115) );
  AND U19115 ( .A(n19349), .B(n17567), .Z(n17651) );
  XNOR U19116 ( .A(n19274), .B(n19113), .Z(n19276) );
  XOR U19117 ( .A(n19277), .B(n19278), .Z(n19113) );
  IV U19118 ( .A(n19279), .Z(n19278) );
  XOR U19119 ( .A(n19280), .B(n19281), .Z(n19274) );
  ANDN U19120 ( .A(n19282), .B(n19121), .Z(n19281) );
  XNOR U19121 ( .A(n19280), .B(n17765), .Z(n19121) );
  AND U19122 ( .A(n19349), .B(n17688), .Z(n17765) );
  XNOR U19123 ( .A(n19280), .B(n19119), .Z(n19282) );
  XOR U19124 ( .A(n19283), .B(n19284), .Z(n19119) );
  IV U19125 ( .A(n19285), .Z(n19284) );
  XOR U19126 ( .A(n19286), .B(n19287), .Z(n19280) );
  ANDN U19127 ( .A(n19288), .B(n19127), .Z(n19287) );
  XNOR U19128 ( .A(n19286), .B(n17884), .Z(n19127) );
  AND U19129 ( .A(n19349), .B(n17814), .Z(n17884) );
  XNOR U19130 ( .A(n19286), .B(n19125), .Z(n19288) );
  XOR U19131 ( .A(n19289), .B(n19290), .Z(n19125) );
  IV U19132 ( .A(n19291), .Z(n19290) );
  XOR U19133 ( .A(n19292), .B(n19293), .Z(n19286) );
  ANDN U19134 ( .A(n19294), .B(n19133), .Z(n19293) );
  XNOR U19135 ( .A(n19292), .B(n18008), .Z(n19133) );
  AND U19136 ( .A(n19349), .B(n17945), .Z(n18008) );
  XNOR U19137 ( .A(n19292), .B(n19131), .Z(n19294) );
  XOR U19138 ( .A(n19295), .B(n19296), .Z(n19131) );
  IV U19139 ( .A(n19297), .Z(n19296) );
  XOR U19140 ( .A(n19298), .B(n19299), .Z(n19292) );
  ANDN U19141 ( .A(n19300), .B(n19139), .Z(n19299) );
  XNOR U19142 ( .A(n19298), .B(n18137), .Z(n19139) );
  AND U19143 ( .A(n19349), .B(n18081), .Z(n18137) );
  XNOR U19144 ( .A(n19298), .B(n19137), .Z(n19300) );
  XOR U19145 ( .A(n19301), .B(n19302), .Z(n19137) );
  IV U19146 ( .A(n19303), .Z(n19302) );
  XOR U19147 ( .A(n19304), .B(n19305), .Z(n19298) );
  ANDN U19148 ( .A(n19306), .B(n19145), .Z(n19305) );
  XNOR U19149 ( .A(n19304), .B(n18271), .Z(n19145) );
  AND U19150 ( .A(n19349), .B(n18222), .Z(n18271) );
  XNOR U19151 ( .A(n19304), .B(n19143), .Z(n19306) );
  XOR U19152 ( .A(n19307), .B(n19308), .Z(n19143) );
  IV U19153 ( .A(n19309), .Z(n19308) );
  XOR U19154 ( .A(n19310), .B(n19311), .Z(n19304) );
  ANDN U19155 ( .A(n19312), .B(n19151), .Z(n19311) );
  XNOR U19156 ( .A(n19310), .B(n18410), .Z(n19151) );
  AND U19157 ( .A(n19349), .B(n18368), .Z(n18410) );
  XNOR U19158 ( .A(n19310), .B(n19149), .Z(n19312) );
  XOR U19159 ( .A(n19313), .B(n19314), .Z(n19149) );
  IV U19160 ( .A(n19315), .Z(n19314) );
  XOR U19161 ( .A(n19316), .B(n19317), .Z(n19310) );
  ANDN U19162 ( .A(n19318), .B(n19157), .Z(n19317) );
  XNOR U19163 ( .A(n19316), .B(n18554), .Z(n19157) );
  AND U19164 ( .A(n19349), .B(n18519), .Z(n18554) );
  XNOR U19165 ( .A(n19316), .B(n19155), .Z(n19318) );
  XOR U19166 ( .A(n19319), .B(n19320), .Z(n19155) );
  IV U19167 ( .A(n19321), .Z(n19320) );
  XOR U19168 ( .A(n19322), .B(n19323), .Z(n19316) );
  ANDN U19169 ( .A(n19324), .B(n19163), .Z(n19323) );
  XNOR U19170 ( .A(n19322), .B(n18703), .Z(n19163) );
  AND U19171 ( .A(n19349), .B(n18675), .Z(n18703) );
  XNOR U19172 ( .A(n19322), .B(n19161), .Z(n19324) );
  XOR U19173 ( .A(n19325), .B(n19326), .Z(n19161) );
  IV U19174 ( .A(n19327), .Z(n19326) );
  XOR U19175 ( .A(n19328), .B(n19329), .Z(n19322) );
  ANDN U19176 ( .A(n19330), .B(n19169), .Z(n19329) );
  XNOR U19177 ( .A(n19328), .B(n18857), .Z(n19169) );
  AND U19178 ( .A(n19349), .B(n18836), .Z(n18857) );
  XNOR U19179 ( .A(n19328), .B(n19167), .Z(n19330) );
  XOR U19180 ( .A(n19331), .B(n19332), .Z(n19167) );
  IV U19181 ( .A(n19333), .Z(n19332) );
  XOR U19182 ( .A(n19334), .B(n19335), .Z(n19328) );
  ANDN U19183 ( .A(n19336), .B(n19176), .Z(n19335) );
  XNOR U19184 ( .A(n19334), .B(n19016), .Z(n19176) );
  AND U19185 ( .A(n19349), .B(n19002), .Z(n19016) );
  XNOR U19186 ( .A(n19334), .B(n19174), .Z(n19336) );
  XOR U19187 ( .A(n19337), .B(n19338), .Z(n19174) );
  IV U19188 ( .A(n19339), .Z(n19338) );
  XOR U19189 ( .A(n19340), .B(n19341), .Z(n19334) );
  ANDN U19190 ( .A(n19342), .B(n19183), .Z(n19341) );
  XNOR U19191 ( .A(n19340), .B(n19180), .Z(n19183) );
  AND U19192 ( .A(n19349), .B(n19173), .Z(n19180) );
  XNOR U19193 ( .A(n19340), .B(n19181), .Z(n19342) );
  XOR U19194 ( .A(n19343), .B(n19344), .Z(n19181) );
  IV U19195 ( .A(n19345), .Z(n19344) );
  XOR U19196 ( .A(n19346), .B(n19347), .Z(n19340) );
  ANDN U19197 ( .A(n19348), .B(n19190), .Z(n19347) );
  XNOR U19198 ( .A(n19346), .B(n19349), .Z(n19190) );
  XNOR U19199 ( .A(n19346), .B(n19188), .Z(n19348) );
  XOR U19200 ( .A(n19350), .B(n19351), .Z(n19188) );
  IV U19201 ( .A(n19352), .Z(n19351) );
  XOR U19202 ( .A(n19353), .B(n19354), .Z(n19346) );
  ANDN U19203 ( .A(n19355), .B(n19196), .Z(n19354) );
  XNOR U19204 ( .A(n19353), .B(n19356), .Z(n19196) );
  XNOR U19205 ( .A(n19353), .B(n19194), .Z(n19355) );
  XOR U19206 ( .A(n19357), .B(n19358), .Z(n19194) );
  IV U19207 ( .A(n19359), .Z(n19358) );
  XOR U19208 ( .A(n19360), .B(n19361), .Z(n19353) );
  NANDN U19209 ( .B(n19200), .A(n19362), .Z(n19360) );
  XOR U19210 ( .A(n19361), .B(n19198), .Z(n19362) );
  XOR U19211 ( .A(n19363), .B(n19364), .Z(n19198) );
  IV U19212 ( .A(n19365), .Z(n19364) );
  XNOR U19213 ( .A(n19366), .B(n19361), .Z(n19200) );
  OR U19214 ( .A(n13247), .B(n13248), .Z(n19361) );
  XOR U19215 ( .A(n19367), .B(n19368), .Z(n13247) );
  IV U19216 ( .A(n19369), .Z(n19368) );
  NAND U19217 ( .A(n16747), .B(n19349), .Z(n19366) );
  XOR U19218 ( .A(n16745), .B(n19370), .Z(n16740) );
  IV U19219 ( .A(n16744), .Z(n19370) );
  XNOR U19220 ( .A(n16741), .B(n16759), .Z(n16744) );
  AND U19221 ( .A(n19478), .B(n13553), .Z(n16759) );
  XOR U19222 ( .A(n19371), .B(n19372), .Z(n16741) );
  ANDN U19223 ( .A(n19373), .B(n19207), .Z(n19372) );
  XNOR U19224 ( .A(n19371), .B(n16775), .Z(n19207) );
  AND U19225 ( .A(n19478), .B(n13636), .Z(n16775) );
  XNOR U19226 ( .A(n19371), .B(n19205), .Z(n19373) );
  XNOR U19227 ( .A(n19374), .B(n9724), .Z(n19205) );
  XOR U19228 ( .A(n19375), .B(n19376), .Z(n19371) );
  ANDN U19229 ( .A(n19377), .B(n19213), .Z(n19376) );
  XNOR U19230 ( .A(n19375), .B(n16801), .Z(n19213) );
  AND U19231 ( .A(n19478), .B(n13745), .Z(n16801) );
  XNOR U19232 ( .A(n19375), .B(n19211), .Z(n19377) );
  XNOR U19233 ( .A(n19378), .B(n9922), .Z(n19211) );
  XOR U19234 ( .A(n19379), .B(n19380), .Z(n19375) );
  ANDN U19235 ( .A(n19381), .B(n19219), .Z(n19380) );
  XNOR U19236 ( .A(n19379), .B(n16834), .Z(n19219) );
  AND U19237 ( .A(n19478), .B(n13880), .Z(n16834) );
  XNOR U19238 ( .A(n19379), .B(n19217), .Z(n19381) );
  XNOR U19239 ( .A(n19382), .B(n10114), .Z(n19217) );
  XOR U19240 ( .A(n19383), .B(n19384), .Z(n19379) );
  ANDN U19241 ( .A(n19385), .B(n19225), .Z(n19384) );
  XNOR U19242 ( .A(n19383), .B(n16874), .Z(n19225) );
  AND U19243 ( .A(n19478), .B(n14041), .Z(n16874) );
  XNOR U19244 ( .A(n19383), .B(n19223), .Z(n19385) );
  XNOR U19245 ( .A(n19386), .B(n10299), .Z(n19223) );
  XOR U19246 ( .A(n19387), .B(n19388), .Z(n19383) );
  ANDN U19247 ( .A(n19389), .B(n19231), .Z(n19388) );
  XNOR U19248 ( .A(n19387), .B(n16921), .Z(n19231) );
  AND U19249 ( .A(n19478), .B(n14228), .Z(n16921) );
  XNOR U19250 ( .A(n19387), .B(n19229), .Z(n19389) );
  XNOR U19251 ( .A(n19390), .B(n10478), .Z(n19229) );
  XOR U19252 ( .A(n19391), .B(n19392), .Z(n19387) );
  ANDN U19253 ( .A(n19393), .B(n19237), .Z(n19392) );
  XNOR U19254 ( .A(n19391), .B(n16975), .Z(n19237) );
  AND U19255 ( .A(n19478), .B(n14441), .Z(n16975) );
  XNOR U19256 ( .A(n19391), .B(n19235), .Z(n19393) );
  XNOR U19257 ( .A(n19394), .B(n10650), .Z(n19235) );
  XOR U19258 ( .A(n19395), .B(n19396), .Z(n19391) );
  ANDN U19259 ( .A(n19397), .B(n19243), .Z(n19396) );
  XNOR U19260 ( .A(n19395), .B(n17036), .Z(n19243) );
  AND U19261 ( .A(n19478), .B(n14680), .Z(n17036) );
  XNOR U19262 ( .A(n19395), .B(n19241), .Z(n19397) );
  XNOR U19263 ( .A(n19398), .B(n10816), .Z(n19241) );
  XOR U19264 ( .A(n19399), .B(n19400), .Z(n19395) );
  ANDN U19265 ( .A(n19401), .B(n19249), .Z(n19400) );
  XNOR U19266 ( .A(n19399), .B(n17104), .Z(n19249) );
  AND U19267 ( .A(n19478), .B(n14945), .Z(n17104) );
  XNOR U19268 ( .A(n19399), .B(n19247), .Z(n19401) );
  XNOR U19269 ( .A(n19402), .B(n10975), .Z(n19247) );
  XOR U19270 ( .A(n19403), .B(n19404), .Z(n19399) );
  ANDN U19271 ( .A(n19405), .B(n19255), .Z(n19404) );
  XNOR U19272 ( .A(n19403), .B(n17179), .Z(n19255) );
  AND U19273 ( .A(n19478), .B(n15236), .Z(n17179) );
  XNOR U19274 ( .A(n19403), .B(n19253), .Z(n19405) );
  XNOR U19275 ( .A(n19406), .B(n11128), .Z(n19253) );
  XOR U19276 ( .A(n19407), .B(n19408), .Z(n19403) );
  ANDN U19277 ( .A(n19409), .B(n19261), .Z(n19408) );
  XNOR U19278 ( .A(n19407), .B(n17261), .Z(n19261) );
  AND U19279 ( .A(n19478), .B(n15553), .Z(n17261) );
  XNOR U19280 ( .A(n19407), .B(n19259), .Z(n19409) );
  XNOR U19281 ( .A(n19410), .B(n11274), .Z(n19259) );
  XOR U19282 ( .A(n19411), .B(n19412), .Z(n19407) );
  ANDN U19283 ( .A(n19413), .B(n19267), .Z(n19412) );
  XNOR U19284 ( .A(n19411), .B(n17350), .Z(n19267) );
  AND U19285 ( .A(n19478), .B(n15896), .Z(n17350) );
  XNOR U19286 ( .A(n19411), .B(n19265), .Z(n19413) );
  XNOR U19287 ( .A(n19414), .B(n11414), .Z(n19265) );
  XOR U19288 ( .A(n19415), .B(n19416), .Z(n19411) );
  ANDN U19289 ( .A(n19417), .B(n19273), .Z(n19416) );
  XNOR U19290 ( .A(n19415), .B(n17446), .Z(n19273) );
  AND U19291 ( .A(n19478), .B(n16265), .Z(n17446) );
  XNOR U19292 ( .A(n19415), .B(n19271), .Z(n19417) );
  XNOR U19293 ( .A(n19418), .B(n11547), .Z(n19271) );
  XOR U19294 ( .A(n19419), .B(n19420), .Z(n19415) );
  ANDN U19295 ( .A(n19421), .B(n19279), .Z(n19420) );
  XNOR U19296 ( .A(n19419), .B(n17549), .Z(n19279) );
  AND U19297 ( .A(n19478), .B(n16657), .Z(n17549) );
  XNOR U19298 ( .A(n19419), .B(n19277), .Z(n19421) );
  XNOR U19299 ( .A(n19422), .B(n11674), .Z(n19277) );
  XOR U19300 ( .A(n19423), .B(n19424), .Z(n19419) );
  ANDN U19301 ( .A(n19425), .B(n19285), .Z(n19424) );
  XNOR U19302 ( .A(n19423), .B(n17658), .Z(n19285) );
  AND U19303 ( .A(n19478), .B(n17567), .Z(n17658) );
  XNOR U19304 ( .A(n19423), .B(n19283), .Z(n19425) );
  XNOR U19305 ( .A(n19426), .B(n11687), .Z(n19283) );
  XOR U19306 ( .A(n19427), .B(n19428), .Z(n19423) );
  ANDN U19307 ( .A(n19429), .B(n19291), .Z(n19428) );
  XNOR U19308 ( .A(n19427), .B(n17772), .Z(n19291) );
  AND U19309 ( .A(n19478), .B(n17688), .Z(n17772) );
  XNOR U19310 ( .A(n19427), .B(n19289), .Z(n19429) );
  XNOR U19311 ( .A(n19430), .B(n11820), .Z(n19289) );
  XOR U19312 ( .A(n19431), .B(n19432), .Z(n19427) );
  ANDN U19313 ( .A(n19433), .B(n19297), .Z(n19432) );
  XNOR U19314 ( .A(n19431), .B(n17891), .Z(n19297) );
  AND U19315 ( .A(n19478), .B(n17814), .Z(n17891) );
  XNOR U19316 ( .A(n19431), .B(n19295), .Z(n19433) );
  XNOR U19317 ( .A(n19434), .B(n11953), .Z(n19295) );
  XOR U19318 ( .A(n19435), .B(n19436), .Z(n19431) );
  ANDN U19319 ( .A(n19437), .B(n19303), .Z(n19436) );
  XNOR U19320 ( .A(n19435), .B(n18015), .Z(n19303) );
  AND U19321 ( .A(n19478), .B(n17945), .Z(n18015) );
  XNOR U19322 ( .A(n19435), .B(n19301), .Z(n19437) );
  XNOR U19323 ( .A(n19438), .B(n12086), .Z(n19301) );
  XOR U19324 ( .A(n19439), .B(n19440), .Z(n19435) );
  ANDN U19325 ( .A(n19441), .B(n19309), .Z(n19440) );
  XNOR U19326 ( .A(n19439), .B(n18144), .Z(n19309) );
  AND U19327 ( .A(n19478), .B(n18081), .Z(n18144) );
  XNOR U19328 ( .A(n19439), .B(n19307), .Z(n19441) );
  XNOR U19329 ( .A(n19442), .B(n12219), .Z(n19307) );
  XOR U19330 ( .A(n19443), .B(n19444), .Z(n19439) );
  ANDN U19331 ( .A(n19445), .B(n19315), .Z(n19444) );
  XNOR U19332 ( .A(n19443), .B(n18278), .Z(n19315) );
  AND U19333 ( .A(n19478), .B(n18222), .Z(n18278) );
  XNOR U19334 ( .A(n19443), .B(n19313), .Z(n19445) );
  XNOR U19335 ( .A(n19446), .B(n12352), .Z(n19313) );
  XOR U19336 ( .A(n19447), .B(n19448), .Z(n19443) );
  ANDN U19337 ( .A(n19449), .B(n19321), .Z(n19448) );
  XNOR U19338 ( .A(n19447), .B(n18417), .Z(n19321) );
  AND U19339 ( .A(n19478), .B(n18368), .Z(n18417) );
  XNOR U19340 ( .A(n19447), .B(n19319), .Z(n19449) );
  XNOR U19341 ( .A(n19450), .B(n12485), .Z(n19319) );
  XOR U19342 ( .A(n19451), .B(n19452), .Z(n19447) );
  ANDN U19343 ( .A(n19453), .B(n19327), .Z(n19452) );
  XNOR U19344 ( .A(n19451), .B(n18561), .Z(n19327) );
  AND U19345 ( .A(n19478), .B(n18519), .Z(n18561) );
  XNOR U19346 ( .A(n19451), .B(n19325), .Z(n19453) );
  XNOR U19347 ( .A(n19454), .B(n12616), .Z(n19325) );
  XOR U19348 ( .A(n19455), .B(n19456), .Z(n19451) );
  ANDN U19349 ( .A(n19457), .B(n19333), .Z(n19456) );
  XNOR U19350 ( .A(n19455), .B(n18710), .Z(n19333) );
  AND U19351 ( .A(n19478), .B(n18675), .Z(n18710) );
  XNOR U19352 ( .A(n19455), .B(n19331), .Z(n19457) );
  XNOR U19353 ( .A(n19458), .B(n12740), .Z(n19331) );
  XOR U19354 ( .A(n19459), .B(n19460), .Z(n19455) );
  ANDN U19355 ( .A(n19461), .B(n19339), .Z(n19460) );
  XNOR U19356 ( .A(n19459), .B(n18864), .Z(n19339) );
  AND U19357 ( .A(n19478), .B(n18836), .Z(n18864) );
  XNOR U19358 ( .A(n19459), .B(n19337), .Z(n19461) );
  XNOR U19359 ( .A(n19462), .B(n12859), .Z(n19337) );
  XOR U19360 ( .A(n19463), .B(n19464), .Z(n19459) );
  ANDN U19361 ( .A(n19465), .B(n19345), .Z(n19464) );
  XNOR U19362 ( .A(n19463), .B(n19023), .Z(n19345) );
  AND U19363 ( .A(n19478), .B(n19002), .Z(n19023) );
  XNOR U19364 ( .A(n19463), .B(n19343), .Z(n19465) );
  XNOR U19365 ( .A(n19466), .B(n12964), .Z(n19343) );
  XOR U19366 ( .A(n19467), .B(n19468), .Z(n19463) );
  ANDN U19367 ( .A(n19469), .B(n19352), .Z(n19468) );
  XNOR U19368 ( .A(n19467), .B(n19187), .Z(n19352) );
  AND U19369 ( .A(n19478), .B(n19173), .Z(n19187) );
  XNOR U19370 ( .A(n19467), .B(n19350), .Z(n19469) );
  XNOR U19371 ( .A(n19470), .B(n13056), .Z(n19350) );
  XOR U19372 ( .A(n19471), .B(n19472), .Z(n19467) );
  ANDN U19373 ( .A(n19473), .B(n19359), .Z(n19472) );
  XNOR U19374 ( .A(n19471), .B(n19356), .Z(n19359) );
  AND U19375 ( .A(n19478), .B(n19349), .Z(n19356) );
  XNOR U19376 ( .A(n19471), .B(n19357), .Z(n19473) );
  XNOR U19377 ( .A(n19474), .B(n13135), .Z(n19357) );
  XOR U19378 ( .A(n19475), .B(n19476), .Z(n19471) );
  ANDN U19379 ( .A(n19477), .B(n19365), .Z(n19476) );
  XNOR U19380 ( .A(n19475), .B(n19478), .Z(n19365) );
  XNOR U19381 ( .A(n19475), .B(n19363), .Z(n19477) );
  XNOR U19382 ( .A(n19479), .B(n13200), .Z(n19363) );
  XNOR U19383 ( .A(n19480), .B(n19481), .Z(n19475) );
  NANDN U19384 ( .B(n19369), .A(n19482), .Z(n19480) );
  XNOR U19385 ( .A(n19481), .B(n19367), .Z(n19482) );
  XNOR U19386 ( .A(n19483), .B(n13248), .Z(n19367) );
  XOR U19387 ( .A(n19484), .B(n19481), .Z(n19369) );
  NOR U19388 ( .A(n13288), .B(n13287), .Z(n19481) );
  XOR U19389 ( .A(n19485), .B(n13287), .Z(n13288) );
  IV U19390 ( .A(n19486), .Z(n19485) );
  NAND U19391 ( .A(n16747), .B(n19478), .Z(n19484) );
  XNOR U19392 ( .A(n16751), .B(n9519), .Z(n16745) );
  NANDN U19393 ( .B(n13320), .A(n13470), .Z(n9519) );
  XNOR U19394 ( .A(n16748), .B(n19487), .Z(n16751) );
  AND U19395 ( .A(n13496), .B(n16747), .Z(n19487) );
  XOR U19396 ( .A(n19488), .B(n19489), .Z(n16748) );
  ANDN U19397 ( .A(n19490), .B(n19374), .Z(n19489) );
  XNOR U19398 ( .A(n19488), .B(n19491), .Z(n19374) );
  AND U19399 ( .A(n13553), .B(n16747), .Z(n19491) );
  XNOR U19400 ( .A(n9724), .B(n19488), .Z(n19490) );
  NANDN U19401 ( .B(n13320), .A(n13496), .Z(n9724) );
  XOR U19402 ( .A(n19492), .B(n19493), .Z(n13496) );
  ANDN U19403 ( .A(n19494), .B(n19495), .Z(n19493) );
  XNOR U19404 ( .A(n19492), .B(n19496), .Z(n19494) );
  XOR U19405 ( .A(n19497), .B(n19498), .Z(n19488) );
  ANDN U19406 ( .A(n19499), .B(n19378), .Z(n19498) );
  XNOR U19407 ( .A(n19497), .B(n19500), .Z(n19378) );
  AND U19408 ( .A(n13636), .B(n16747), .Z(n19500) );
  XNOR U19409 ( .A(n9922), .B(n19497), .Z(n19499) );
  NANDN U19410 ( .B(n13320), .A(n13553), .Z(n9922) );
  XOR U19411 ( .A(n19501), .B(n19502), .Z(n13553) );
  ANDN U19412 ( .A(n19503), .B(n19495), .Z(n19502) );
  XNOR U19413 ( .A(n19501), .B(n19504), .Z(n19503) );
  XOR U19414 ( .A(n19505), .B(n19506), .Z(n19497) );
  ANDN U19415 ( .A(n19507), .B(n19382), .Z(n19506) );
  XNOR U19416 ( .A(n19505), .B(n19508), .Z(n19382) );
  AND U19417 ( .A(n13745), .B(n16747), .Z(n19508) );
  XNOR U19418 ( .A(n10114), .B(n19505), .Z(n19507) );
  NANDN U19419 ( .B(n13320), .A(n13636), .Z(n10114) );
  XOR U19420 ( .A(n19509), .B(n19510), .Z(n13636) );
  ANDN U19421 ( .A(n19511), .B(n19495), .Z(n19510) );
  XNOR U19422 ( .A(n19509), .B(n19512), .Z(n19511) );
  XOR U19423 ( .A(n19513), .B(n19514), .Z(n19505) );
  ANDN U19424 ( .A(n19515), .B(n19386), .Z(n19514) );
  XNOR U19425 ( .A(n19513), .B(n19516), .Z(n19386) );
  AND U19426 ( .A(n13880), .B(n16747), .Z(n19516) );
  XNOR U19427 ( .A(n10299), .B(n19513), .Z(n19515) );
  NANDN U19428 ( .B(n13320), .A(n13745), .Z(n10299) );
  XOR U19429 ( .A(n19517), .B(n19518), .Z(n13745) );
  ANDN U19430 ( .A(n19519), .B(n19495), .Z(n19518) );
  XNOR U19431 ( .A(n19517), .B(n19520), .Z(n19519) );
  XOR U19432 ( .A(n19521), .B(n19522), .Z(n19513) );
  ANDN U19433 ( .A(n19523), .B(n19390), .Z(n19522) );
  XNOR U19434 ( .A(n19521), .B(n19524), .Z(n19390) );
  AND U19435 ( .A(n14041), .B(n16747), .Z(n19524) );
  XNOR U19436 ( .A(n10478), .B(n19521), .Z(n19523) );
  NANDN U19437 ( .B(n13320), .A(n13880), .Z(n10478) );
  XOR U19438 ( .A(n19525), .B(n19526), .Z(n13880) );
  ANDN U19439 ( .A(n19527), .B(n19495), .Z(n19526) );
  XNOR U19440 ( .A(n19525), .B(n19528), .Z(n19527) );
  XOR U19441 ( .A(n19529), .B(n19530), .Z(n19521) );
  ANDN U19442 ( .A(n19531), .B(n19394), .Z(n19530) );
  XNOR U19443 ( .A(n19529), .B(n19532), .Z(n19394) );
  AND U19444 ( .A(n14228), .B(n16747), .Z(n19532) );
  XNOR U19445 ( .A(n10650), .B(n19529), .Z(n19531) );
  NANDN U19446 ( .B(n13320), .A(n14041), .Z(n10650) );
  XOR U19447 ( .A(n19533), .B(n19534), .Z(n14041) );
  ANDN U19448 ( .A(n19535), .B(n19495), .Z(n19534) );
  XNOR U19449 ( .A(n19533), .B(n19536), .Z(n19535) );
  XOR U19450 ( .A(n19537), .B(n19538), .Z(n19529) );
  ANDN U19451 ( .A(n19539), .B(n19398), .Z(n19538) );
  XNOR U19452 ( .A(n19537), .B(n19540), .Z(n19398) );
  AND U19453 ( .A(n14441), .B(n16747), .Z(n19540) );
  XNOR U19454 ( .A(n10816), .B(n19537), .Z(n19539) );
  NANDN U19455 ( .B(n13320), .A(n14228), .Z(n10816) );
  XOR U19456 ( .A(n19541), .B(n19542), .Z(n14228) );
  ANDN U19457 ( .A(n19543), .B(n19495), .Z(n19542) );
  XNOR U19458 ( .A(n19541), .B(n19544), .Z(n19543) );
  XOR U19459 ( .A(n19545), .B(n19546), .Z(n19537) );
  ANDN U19460 ( .A(n19547), .B(n19402), .Z(n19546) );
  XNOR U19461 ( .A(n19545), .B(n19548), .Z(n19402) );
  AND U19462 ( .A(n14680), .B(n16747), .Z(n19548) );
  XNOR U19463 ( .A(n10975), .B(n19545), .Z(n19547) );
  NANDN U19464 ( .B(n13320), .A(n14441), .Z(n10975) );
  XOR U19465 ( .A(n19549), .B(n19550), .Z(n14441) );
  ANDN U19466 ( .A(n19551), .B(n19495), .Z(n19550) );
  XNOR U19467 ( .A(n19549), .B(n19552), .Z(n19551) );
  XOR U19468 ( .A(n19553), .B(n19554), .Z(n19545) );
  ANDN U19469 ( .A(n19555), .B(n19406), .Z(n19554) );
  XNOR U19470 ( .A(n19553), .B(n19556), .Z(n19406) );
  AND U19471 ( .A(n14945), .B(n16747), .Z(n19556) );
  XNOR U19472 ( .A(n11128), .B(n19553), .Z(n19555) );
  NANDN U19473 ( .B(n13320), .A(n14680), .Z(n11128) );
  XOR U19474 ( .A(n19557), .B(n19558), .Z(n14680) );
  ANDN U19475 ( .A(n19559), .B(n19495), .Z(n19558) );
  XNOR U19476 ( .A(n19557), .B(n19560), .Z(n19559) );
  XOR U19477 ( .A(n19561), .B(n19562), .Z(n19553) );
  ANDN U19478 ( .A(n19563), .B(n19410), .Z(n19562) );
  XNOR U19479 ( .A(n19561), .B(n19564), .Z(n19410) );
  AND U19480 ( .A(n15236), .B(n16747), .Z(n19564) );
  XNOR U19481 ( .A(n11274), .B(n19561), .Z(n19563) );
  NANDN U19482 ( .B(n13320), .A(n14945), .Z(n11274) );
  XOR U19483 ( .A(n19565), .B(n19566), .Z(n14945) );
  ANDN U19484 ( .A(n19567), .B(n19495), .Z(n19566) );
  XNOR U19485 ( .A(n19565), .B(n19568), .Z(n19567) );
  XOR U19486 ( .A(n19569), .B(n19570), .Z(n19561) );
  ANDN U19487 ( .A(n19571), .B(n19414), .Z(n19570) );
  XNOR U19488 ( .A(n19569), .B(n19572), .Z(n19414) );
  AND U19489 ( .A(n15553), .B(n16747), .Z(n19572) );
  XNOR U19490 ( .A(n11414), .B(n19569), .Z(n19571) );
  NANDN U19491 ( .B(n13320), .A(n15236), .Z(n11414) );
  XOR U19492 ( .A(n19573), .B(n19574), .Z(n15236) );
  ANDN U19493 ( .A(n19575), .B(n19495), .Z(n19574) );
  XNOR U19494 ( .A(n19573), .B(n19576), .Z(n19575) );
  XOR U19495 ( .A(n19577), .B(n19578), .Z(n19569) );
  ANDN U19496 ( .A(n19579), .B(n19418), .Z(n19578) );
  XNOR U19497 ( .A(n19577), .B(n19580), .Z(n19418) );
  AND U19498 ( .A(n15896), .B(n16747), .Z(n19580) );
  XNOR U19499 ( .A(n11547), .B(n19577), .Z(n19579) );
  NANDN U19500 ( .B(n13320), .A(n15553), .Z(n11547) );
  XOR U19501 ( .A(n19581), .B(n19582), .Z(n15553) );
  ANDN U19502 ( .A(n19583), .B(n19495), .Z(n19582) );
  XNOR U19503 ( .A(n19581), .B(n19584), .Z(n19583) );
  XOR U19504 ( .A(n19585), .B(n19586), .Z(n19577) );
  ANDN U19505 ( .A(n19587), .B(n19422), .Z(n19586) );
  XNOR U19506 ( .A(n19585), .B(n19588), .Z(n19422) );
  AND U19507 ( .A(n16265), .B(n16747), .Z(n19588) );
  XNOR U19508 ( .A(n11674), .B(n19585), .Z(n19587) );
  NANDN U19509 ( .B(n13320), .A(n15896), .Z(n11674) );
  XOR U19510 ( .A(n19589), .B(n19590), .Z(n15896) );
  ANDN U19511 ( .A(n19591), .B(n19495), .Z(n19590) );
  XNOR U19512 ( .A(n19589), .B(n19592), .Z(n19591) );
  XOR U19513 ( .A(n19593), .B(n19594), .Z(n19585) );
  ANDN U19514 ( .A(n19595), .B(n19426), .Z(n19594) );
  XNOR U19515 ( .A(n19593), .B(n19596), .Z(n19426) );
  AND U19516 ( .A(n16657), .B(n16747), .Z(n19596) );
  XNOR U19517 ( .A(n11687), .B(n19593), .Z(n19595) );
  NANDN U19518 ( .B(n13320), .A(n16265), .Z(n11687) );
  XOR U19519 ( .A(n19597), .B(n19598), .Z(n16265) );
  ANDN U19520 ( .A(n19599), .B(n19495), .Z(n19598) );
  XNOR U19521 ( .A(n19597), .B(n19600), .Z(n19599) );
  XOR U19522 ( .A(n19601), .B(n19602), .Z(n19593) );
  ANDN U19523 ( .A(n19603), .B(n19430), .Z(n19602) );
  XNOR U19524 ( .A(n19601), .B(n19604), .Z(n19430) );
  AND U19525 ( .A(n17567), .B(n16747), .Z(n19604) );
  XNOR U19526 ( .A(n11820), .B(n19601), .Z(n19603) );
  NANDN U19527 ( .B(n13320), .A(n16657), .Z(n11820) );
  XOR U19528 ( .A(n19605), .B(n19606), .Z(n16657) );
  ANDN U19529 ( .A(n19607), .B(n19495), .Z(n19606) );
  XNOR U19530 ( .A(n19605), .B(n19608), .Z(n19607) );
  XOR U19531 ( .A(n19609), .B(n19610), .Z(n19601) );
  ANDN U19532 ( .A(n19611), .B(n19434), .Z(n19610) );
  XNOR U19533 ( .A(n19609), .B(n19612), .Z(n19434) );
  AND U19534 ( .A(n17688), .B(n16747), .Z(n19612) );
  XNOR U19535 ( .A(n11953), .B(n19609), .Z(n19611) );
  NANDN U19536 ( .B(n13320), .A(n17567), .Z(n11953) );
  XOR U19537 ( .A(n19613), .B(n19614), .Z(n17567) );
  ANDN U19538 ( .A(n19615), .B(n19495), .Z(n19614) );
  XNOR U19539 ( .A(n19613), .B(n19616), .Z(n19615) );
  XOR U19540 ( .A(n19617), .B(n19618), .Z(n19609) );
  ANDN U19541 ( .A(n19619), .B(n19438), .Z(n19618) );
  XNOR U19542 ( .A(n19617), .B(n19620), .Z(n19438) );
  AND U19543 ( .A(n17814), .B(n16747), .Z(n19620) );
  XNOR U19544 ( .A(n12086), .B(n19617), .Z(n19619) );
  NANDN U19545 ( .B(n13320), .A(n17688), .Z(n12086) );
  XOR U19546 ( .A(n19621), .B(n19622), .Z(n17688) );
  ANDN U19547 ( .A(n19623), .B(n19495), .Z(n19622) );
  XNOR U19548 ( .A(n19621), .B(n19624), .Z(n19623) );
  XOR U19549 ( .A(n19625), .B(n19626), .Z(n19617) );
  ANDN U19550 ( .A(n19627), .B(n19442), .Z(n19626) );
  XNOR U19551 ( .A(n19625), .B(n19628), .Z(n19442) );
  AND U19552 ( .A(n17945), .B(n16747), .Z(n19628) );
  XNOR U19553 ( .A(n12219), .B(n19625), .Z(n19627) );
  NANDN U19554 ( .B(n13320), .A(n17814), .Z(n12219) );
  XOR U19555 ( .A(n19629), .B(n19630), .Z(n17814) );
  ANDN U19556 ( .A(n19631), .B(n19495), .Z(n19630) );
  XNOR U19557 ( .A(n19629), .B(n19632), .Z(n19631) );
  XOR U19558 ( .A(n19633), .B(n19634), .Z(n19625) );
  ANDN U19559 ( .A(n19635), .B(n19446), .Z(n19634) );
  XNOR U19560 ( .A(n19633), .B(n19636), .Z(n19446) );
  AND U19561 ( .A(n18081), .B(n16747), .Z(n19636) );
  XNOR U19562 ( .A(n12352), .B(n19633), .Z(n19635) );
  NANDN U19563 ( .B(n13320), .A(n17945), .Z(n12352) );
  XOR U19564 ( .A(n19637), .B(n19638), .Z(n17945) );
  ANDN U19565 ( .A(n19639), .B(n19495), .Z(n19638) );
  XNOR U19566 ( .A(n19637), .B(n19640), .Z(n19639) );
  XOR U19567 ( .A(n19641), .B(n19642), .Z(n19633) );
  ANDN U19568 ( .A(n19643), .B(n19450), .Z(n19642) );
  XNOR U19569 ( .A(n19641), .B(n19644), .Z(n19450) );
  AND U19570 ( .A(n18222), .B(n16747), .Z(n19644) );
  XNOR U19571 ( .A(n12485), .B(n19641), .Z(n19643) );
  NANDN U19572 ( .B(n13320), .A(n18081), .Z(n12485) );
  XOR U19573 ( .A(n19645), .B(n19646), .Z(n18081) );
  ANDN U19574 ( .A(n19647), .B(n19495), .Z(n19646) );
  XNOR U19575 ( .A(n19645), .B(n19648), .Z(n19647) );
  XOR U19576 ( .A(n19649), .B(n19650), .Z(n19641) );
  ANDN U19577 ( .A(n19651), .B(n19454), .Z(n19650) );
  XNOR U19578 ( .A(n19649), .B(n19652), .Z(n19454) );
  AND U19579 ( .A(n18368), .B(n16747), .Z(n19652) );
  XNOR U19580 ( .A(n12616), .B(n19649), .Z(n19651) );
  NANDN U19581 ( .B(n13320), .A(n18222), .Z(n12616) );
  XOR U19582 ( .A(n19653), .B(n19654), .Z(n18222) );
  ANDN U19583 ( .A(n19655), .B(n19495), .Z(n19654) );
  XNOR U19584 ( .A(n19653), .B(n19656), .Z(n19655) );
  XOR U19585 ( .A(n19657), .B(n19658), .Z(n19649) );
  ANDN U19586 ( .A(n19659), .B(n19458), .Z(n19658) );
  XNOR U19587 ( .A(n19657), .B(n19660), .Z(n19458) );
  AND U19588 ( .A(n18519), .B(n16747), .Z(n19660) );
  XNOR U19589 ( .A(n12740), .B(n19657), .Z(n19659) );
  NANDN U19590 ( .B(n13320), .A(n18368), .Z(n12740) );
  XOR U19591 ( .A(n19661), .B(n19662), .Z(n18368) );
  ANDN U19592 ( .A(n19663), .B(n19495), .Z(n19662) );
  XNOR U19593 ( .A(n19661), .B(n19664), .Z(n19663) );
  XOR U19594 ( .A(n19665), .B(n19666), .Z(n19657) );
  ANDN U19595 ( .A(n19667), .B(n19462), .Z(n19666) );
  XNOR U19596 ( .A(n19665), .B(n19668), .Z(n19462) );
  AND U19597 ( .A(n18675), .B(n16747), .Z(n19668) );
  XNOR U19598 ( .A(n12859), .B(n19665), .Z(n19667) );
  NANDN U19599 ( .B(n13320), .A(n18519), .Z(n12859) );
  XOR U19600 ( .A(n19669), .B(n19670), .Z(n18519) );
  ANDN U19601 ( .A(n19671), .B(n19495), .Z(n19670) );
  XNOR U19602 ( .A(n19669), .B(n19672), .Z(n19671) );
  XOR U19603 ( .A(n19673), .B(n19674), .Z(n19665) );
  ANDN U19604 ( .A(n19675), .B(n19466), .Z(n19674) );
  XNOR U19605 ( .A(n19673), .B(n19676), .Z(n19466) );
  AND U19606 ( .A(n18836), .B(n16747), .Z(n19676) );
  XNOR U19607 ( .A(n12964), .B(n19673), .Z(n19675) );
  NANDN U19608 ( .B(n13320), .A(n18675), .Z(n12964) );
  XOR U19609 ( .A(n19677), .B(n19678), .Z(n18675) );
  ANDN U19610 ( .A(n19679), .B(n19495), .Z(n19678) );
  XNOR U19611 ( .A(n19677), .B(n19680), .Z(n19679) );
  XOR U19612 ( .A(n19681), .B(n19682), .Z(n19673) );
  ANDN U19613 ( .A(n19683), .B(n19470), .Z(n19682) );
  XNOR U19614 ( .A(n19681), .B(n19684), .Z(n19470) );
  AND U19615 ( .A(n19002), .B(n16747), .Z(n19684) );
  XNOR U19616 ( .A(n13056), .B(n19681), .Z(n19683) );
  NANDN U19617 ( .B(n13320), .A(n18836), .Z(n13056) );
  XOR U19618 ( .A(n19685), .B(n19686), .Z(n18836) );
  ANDN U19619 ( .A(n19687), .B(n19495), .Z(n19686) );
  XNOR U19620 ( .A(n19685), .B(n19688), .Z(n19687) );
  XOR U19621 ( .A(n19689), .B(n19690), .Z(n19681) );
  ANDN U19622 ( .A(n19691), .B(n19474), .Z(n19690) );
  XNOR U19623 ( .A(n19689), .B(n19692), .Z(n19474) );
  AND U19624 ( .A(n19173), .B(n16747), .Z(n19692) );
  XNOR U19625 ( .A(n13135), .B(n19689), .Z(n19691) );
  NANDN U19626 ( .B(n13320), .A(n19002), .Z(n13135) );
  XOR U19627 ( .A(n19693), .B(n19694), .Z(n19002) );
  ANDN U19628 ( .A(n19695), .B(n19495), .Z(n19694) );
  XNOR U19629 ( .A(n19693), .B(n19696), .Z(n19695) );
  XOR U19630 ( .A(n19697), .B(n19698), .Z(n19689) );
  ANDN U19631 ( .A(n19699), .B(n19479), .Z(n19698) );
  XNOR U19632 ( .A(n19697), .B(n19700), .Z(n19479) );
  AND U19633 ( .A(n19349), .B(n16747), .Z(n19700) );
  XNOR U19634 ( .A(n13200), .B(n19697), .Z(n19699) );
  NANDN U19635 ( .B(n13320), .A(n19173), .Z(n13200) );
  XOR U19636 ( .A(n19701), .B(n19702), .Z(n19173) );
  ANDN U19637 ( .A(n19703), .B(n19495), .Z(n19702) );
  XNOR U19638 ( .A(n19701), .B(n19704), .Z(n19703) );
  XOR U19639 ( .A(n19705), .B(n19706), .Z(n19697) );
  ANDN U19640 ( .A(n19707), .B(n19483), .Z(n19706) );
  XNOR U19641 ( .A(n19705), .B(n19708), .Z(n19483) );
  AND U19642 ( .A(n19478), .B(n16747), .Z(n19708) );
  XNOR U19643 ( .A(n13248), .B(n19705), .Z(n19707) );
  NANDN U19644 ( .B(n13320), .A(n19349), .Z(n13248) );
  XOR U19645 ( .A(n19709), .B(n19710), .Z(n19349) );
  ANDN U19646 ( .A(n19711), .B(n19495), .Z(n19710) );
  XNOR U19647 ( .A(n19709), .B(n19712), .Z(n19711) );
  XNOR U19648 ( .A(n19713), .B(n19714), .Z(n19705) );
  NANDN U19649 ( .B(n19486), .A(n19715), .Z(n19713) );
  XNOR U19650 ( .A(n13287), .B(n19714), .Z(n19715) );
  NANDN U19651 ( .B(n13320), .A(n19478), .Z(n13287) );
  XOR U19652 ( .A(n19716), .B(n19717), .Z(n19478) );
  ANDN U19653 ( .A(n19718), .B(n19495), .Z(n19717) );
  XNOR U19654 ( .A(n19716), .B(n19719), .Z(n19718) );
  XOR U19655 ( .A(n19720), .B(n19714), .Z(n19486) );
  ANDN U19656 ( .A(n13453), .B(n13454), .Z(n19714) );
  NANDN U19657 ( .B(n13320), .A(n16747), .Z(n13454) );
  ANDN U19658 ( .A(n16747), .B(n13320), .Z(n13453) );
  NAND U19659 ( .A(n16747), .B(n13470), .Z(n16752) );
  XNOR U19660 ( .A(n19495), .B(n19721), .Z(n13470) );
  ANDN U19661 ( .A(n19722), .B(n19495), .Z(n19721) );
  XNOR U19662 ( .A(n19723), .B(n19724), .Z(n19722) );
  ANDN U19663 ( .A(n19724), .B(n19496), .Z(n19723) );
  XOR U19664 ( .A(n19724), .B(n19492), .Z(n19496) );
  XOR U19665 ( .A(n19725), .B(n19726), .Z(n19724) );
  ANDN U19666 ( .A(n19725), .B(n19504), .Z(n19726) );
  XOR U19667 ( .A(n19725), .B(n19501), .Z(n19504) );
  XOR U19668 ( .A(n19727), .B(n19728), .Z(n19501) );
  XOR U19669 ( .A(n19729), .B(n19730), .Z(n19725) );
  ANDN U19670 ( .A(n19729), .B(n19512), .Z(n19730) );
  XOR U19671 ( .A(n19729), .B(n19509), .Z(n19512) );
  XOR U19672 ( .A(n19731), .B(n19728), .Z(n19509) );
  XOR U19673 ( .A(n19732), .B(n19733), .Z(n19729) );
  ANDN U19674 ( .A(n19732), .B(n19520), .Z(n19733) );
  XOR U19675 ( .A(n19732), .B(n19517), .Z(n19520) );
  XOR U19676 ( .A(n19734), .B(n19728), .Z(n19517) );
  XOR U19677 ( .A(n19735), .B(n19736), .Z(n19732) );
  ANDN U19678 ( .A(n19735), .B(n19528), .Z(n19736) );
  XOR U19679 ( .A(n19735), .B(n19525), .Z(n19528) );
  XOR U19680 ( .A(n19737), .B(n19728), .Z(n19525) );
  XOR U19681 ( .A(n19738), .B(n19739), .Z(n19735) );
  ANDN U19682 ( .A(n19738), .B(n19536), .Z(n19739) );
  XOR U19683 ( .A(n19738), .B(n19533), .Z(n19536) );
  XOR U19684 ( .A(n19740), .B(n19728), .Z(n19533) );
  XOR U19685 ( .A(n19741), .B(n19742), .Z(n19738) );
  ANDN U19686 ( .A(n19741), .B(n19544), .Z(n19742) );
  XOR U19687 ( .A(n19741), .B(n19541), .Z(n19544) );
  XOR U19688 ( .A(n19743), .B(n19728), .Z(n19541) );
  XOR U19689 ( .A(n19744), .B(n19745), .Z(n19741) );
  ANDN U19690 ( .A(n19744), .B(n19552), .Z(n19745) );
  XOR U19691 ( .A(n19744), .B(n19549), .Z(n19552) );
  XOR U19692 ( .A(n19746), .B(n19728), .Z(n19549) );
  XOR U19693 ( .A(n19747), .B(n19748), .Z(n19744) );
  ANDN U19694 ( .A(n19747), .B(n19560), .Z(n19748) );
  XOR U19695 ( .A(n19747), .B(n19557), .Z(n19560) );
  XOR U19696 ( .A(n19749), .B(n19728), .Z(n19557) );
  XOR U19697 ( .A(n19750), .B(n19751), .Z(n19747) );
  ANDN U19698 ( .A(n19750), .B(n19568), .Z(n19751) );
  XOR U19699 ( .A(n19750), .B(n19565), .Z(n19568) );
  XOR U19700 ( .A(n19752), .B(n19728), .Z(n19565) );
  XOR U19701 ( .A(n19753), .B(n19754), .Z(n19750) );
  ANDN U19702 ( .A(n19753), .B(n19576), .Z(n19754) );
  XOR U19703 ( .A(n19753), .B(n19573), .Z(n19576) );
  XOR U19704 ( .A(n19755), .B(n19728), .Z(n19573) );
  XOR U19705 ( .A(n19756), .B(n19757), .Z(n19753) );
  ANDN U19706 ( .A(n19756), .B(n19584), .Z(n19757) );
  XOR U19707 ( .A(n19756), .B(n19581), .Z(n19584) );
  XOR U19708 ( .A(n19758), .B(n19728), .Z(n19581) );
  XOR U19709 ( .A(n19759), .B(n19760), .Z(n19756) );
  ANDN U19710 ( .A(n19759), .B(n19592), .Z(n19760) );
  XOR U19711 ( .A(n19759), .B(n19589), .Z(n19592) );
  XOR U19712 ( .A(n19761), .B(n19728), .Z(n19589) );
  XOR U19713 ( .A(n19762), .B(n19763), .Z(n19759) );
  ANDN U19714 ( .A(n19762), .B(n19600), .Z(n19763) );
  XOR U19715 ( .A(n19762), .B(n19597), .Z(n19600) );
  XOR U19716 ( .A(n19764), .B(n19728), .Z(n19597) );
  XOR U19717 ( .A(n19765), .B(n19766), .Z(n19762) );
  ANDN U19718 ( .A(n19765), .B(n19608), .Z(n19766) );
  XOR U19719 ( .A(n19765), .B(n19605), .Z(n19608) );
  XOR U19720 ( .A(n19767), .B(n19728), .Z(n19605) );
  XOR U19721 ( .A(n19768), .B(n19769), .Z(n19765) );
  ANDN U19722 ( .A(n19768), .B(n19616), .Z(n19769) );
  XOR U19723 ( .A(n19768), .B(n19613), .Z(n19616) );
  XOR U19724 ( .A(n19770), .B(n19728), .Z(n19613) );
  XOR U19725 ( .A(n19771), .B(n19772), .Z(n19768) );
  ANDN U19726 ( .A(n19771), .B(n19624), .Z(n19772) );
  XOR U19727 ( .A(n19771), .B(n19621), .Z(n19624) );
  XOR U19728 ( .A(n19773), .B(n19728), .Z(n19621) );
  XOR U19729 ( .A(n19774), .B(n19775), .Z(n19771) );
  ANDN U19730 ( .A(n19774), .B(n19632), .Z(n19775) );
  XOR U19731 ( .A(n19774), .B(n19629), .Z(n19632) );
  XOR U19732 ( .A(n19776), .B(n19728), .Z(n19629) );
  XOR U19733 ( .A(n19777), .B(n19778), .Z(n19774) );
  ANDN U19734 ( .A(n19777), .B(n19640), .Z(n19778) );
  XOR U19735 ( .A(n19777), .B(n19637), .Z(n19640) );
  XOR U19736 ( .A(n19779), .B(n19728), .Z(n19637) );
  XOR U19737 ( .A(n19780), .B(n19781), .Z(n19777) );
  ANDN U19738 ( .A(n19780), .B(n19648), .Z(n19781) );
  XOR U19739 ( .A(n19780), .B(n19645), .Z(n19648) );
  XOR U19740 ( .A(n19782), .B(n19728), .Z(n19645) );
  XOR U19741 ( .A(n19783), .B(n19784), .Z(n19780) );
  ANDN U19742 ( .A(n19783), .B(n19656), .Z(n19784) );
  XOR U19743 ( .A(n19783), .B(n19653), .Z(n19656) );
  XOR U19744 ( .A(n19785), .B(n19728), .Z(n19653) );
  XOR U19745 ( .A(n19786), .B(n19787), .Z(n19783) );
  ANDN U19746 ( .A(n19786), .B(n19664), .Z(n19787) );
  XOR U19747 ( .A(n19786), .B(n19661), .Z(n19664) );
  XOR U19748 ( .A(n19788), .B(n19728), .Z(n19661) );
  XOR U19749 ( .A(n19789), .B(n19790), .Z(n19786) );
  ANDN U19750 ( .A(n19789), .B(n19672), .Z(n19790) );
  XOR U19751 ( .A(n19789), .B(n19669), .Z(n19672) );
  XOR U19752 ( .A(n19791), .B(n19728), .Z(n19669) );
  XOR U19753 ( .A(n19792), .B(n19793), .Z(n19789) );
  ANDN U19754 ( .A(n19792), .B(n19680), .Z(n19793) );
  XOR U19755 ( .A(n19792), .B(n19677), .Z(n19680) );
  XOR U19756 ( .A(n19794), .B(n19728), .Z(n19677) );
  XOR U19757 ( .A(n19795), .B(n19796), .Z(n19792) );
  ANDN U19758 ( .A(n19795), .B(n19688), .Z(n19796) );
  XOR U19759 ( .A(n19795), .B(n19685), .Z(n19688) );
  XNOR U19760 ( .A(n19797), .B(e_input[15]), .Z(n19685) );
  XOR U19761 ( .A(n19798), .B(n19799), .Z(n19795) );
  ANDN U19762 ( .A(n19798), .B(n19696), .Z(n19799) );
  XOR U19763 ( .A(n19798), .B(n19693), .Z(n19696) );
  XNOR U19764 ( .A(n19800), .B(e_input[14]), .Z(n19693) );
  XOR U19765 ( .A(n19801), .B(n19802), .Z(n19798) );
  ANDN U19766 ( .A(n19801), .B(n19704), .Z(n19802) );
  XOR U19767 ( .A(n19801), .B(n19701), .Z(n19704) );
  XNOR U19768 ( .A(n19803), .B(e_input[13]), .Z(n19701) );
  XOR U19769 ( .A(n19804), .B(n19805), .Z(n19801) );
  ANDN U19770 ( .A(n19804), .B(n19712), .Z(n19805) );
  XOR U19771 ( .A(n19804), .B(n19709), .Z(n19712) );
  XNOR U19772 ( .A(n19806), .B(e_input[12]), .Z(n19709) );
  XNOR U19773 ( .A(n19807), .B(n19808), .Z(n19804) );
  NOR U19774 ( .A(n19807), .B(n19719), .Z(n19808) );
  XNOR U19775 ( .A(n19807), .B(n19716), .Z(n19719) );
  XNOR U19776 ( .A(n19809), .B(e_input[11]), .Z(n19716) );
  XNOR U19777 ( .A(n13320), .B(n19810), .Z(n19807) );
  NOR U19778 ( .A(n19811), .B(n19812), .Z(n19810) );
  IV U19779 ( .A(n19811), .Z(n13320) );
  XNOR U19780 ( .A(n19813), .B(n19814), .Z(n16747) );
  ANDN U19781 ( .A(n19815), .B(n19495), .Z(n19814) );
  XOR U19782 ( .A(n19816), .B(n19817), .Z(n19495) );
  AND U19783 ( .A(n19818), .B(n19819), .Z(n19817) );
  XOR U19784 ( .A(n19728), .B(g_input[30]), .Z(n19819) );
  XNOR U19785 ( .A(n19492), .B(n19816), .Z(n19818) );
  XOR U19786 ( .A(n19820), .B(e_input[16]), .Z(n19492) );
  XOR U19787 ( .A(n19821), .B(n19822), .Z(n19816) );
  ANDN U19788 ( .A(n19823), .B(n19820), .Z(n19822) );
  XOR U19789 ( .A(n19821), .B(g_input[30]), .Z(n19820) );
  XNOR U19790 ( .A(n19728), .B(n19821), .Z(n19823) );
  XOR U19791 ( .A(n19824), .B(n19825), .Z(n19821) );
  AND U19792 ( .A(n19727), .B(n19826), .Z(n19825) );
  XNOR U19793 ( .A(n19728), .B(n19824), .Z(n19826) );
  XNOR U19794 ( .A(n19824), .B(g_input[29]), .Z(n19727) );
  XOR U19795 ( .A(n19827), .B(n19828), .Z(n19824) );
  AND U19796 ( .A(n19731), .B(n19829), .Z(n19828) );
  XNOR U19797 ( .A(n19728), .B(n19827), .Z(n19829) );
  XNOR U19798 ( .A(n19827), .B(g_input[28]), .Z(n19731) );
  XOR U19799 ( .A(n19830), .B(n19831), .Z(n19827) );
  AND U19800 ( .A(n19734), .B(n19832), .Z(n19831) );
  XNOR U19801 ( .A(n19728), .B(n19830), .Z(n19832) );
  XNOR U19802 ( .A(n19830), .B(g_input[27]), .Z(n19734) );
  XOR U19803 ( .A(n19833), .B(n19834), .Z(n19830) );
  AND U19804 ( .A(n19737), .B(n19835), .Z(n19834) );
  XNOR U19805 ( .A(n19728), .B(n19833), .Z(n19835) );
  XNOR U19806 ( .A(n19833), .B(g_input[26]), .Z(n19737) );
  XOR U19807 ( .A(n19836), .B(n19837), .Z(n19833) );
  AND U19808 ( .A(n19740), .B(n19838), .Z(n19837) );
  XNOR U19809 ( .A(n19728), .B(n19836), .Z(n19838) );
  XNOR U19810 ( .A(n19836), .B(g_input[25]), .Z(n19740) );
  XOR U19811 ( .A(n19839), .B(n19840), .Z(n19836) );
  AND U19812 ( .A(n19743), .B(n19841), .Z(n19840) );
  XNOR U19813 ( .A(n19728), .B(n19839), .Z(n19841) );
  XNOR U19814 ( .A(n19839), .B(g_input[24]), .Z(n19743) );
  XOR U19815 ( .A(n19842), .B(n19843), .Z(n19839) );
  AND U19816 ( .A(n19746), .B(n19844), .Z(n19843) );
  XNOR U19817 ( .A(n19728), .B(n19842), .Z(n19844) );
  XNOR U19818 ( .A(n19842), .B(g_input[23]), .Z(n19746) );
  XOR U19819 ( .A(n19845), .B(n19846), .Z(n19842) );
  AND U19820 ( .A(n19749), .B(n19847), .Z(n19846) );
  XNOR U19821 ( .A(n19728), .B(n19845), .Z(n19847) );
  XNOR U19822 ( .A(n19845), .B(g_input[22]), .Z(n19749) );
  XOR U19823 ( .A(n19848), .B(n19849), .Z(n19845) );
  AND U19824 ( .A(n19752), .B(n19850), .Z(n19849) );
  XNOR U19825 ( .A(n19728), .B(n19848), .Z(n19850) );
  XNOR U19826 ( .A(n19848), .B(g_input[21]), .Z(n19752) );
  XOR U19827 ( .A(n19851), .B(n19852), .Z(n19848) );
  AND U19828 ( .A(n19755), .B(n19853), .Z(n19852) );
  XNOR U19829 ( .A(n19728), .B(n19851), .Z(n19853) );
  XNOR U19830 ( .A(n19851), .B(g_input[20]), .Z(n19755) );
  XOR U19831 ( .A(n19854), .B(n19855), .Z(n19851) );
  AND U19832 ( .A(n19758), .B(n19856), .Z(n19855) );
  XNOR U19833 ( .A(n19728), .B(n19854), .Z(n19856) );
  XNOR U19834 ( .A(n19854), .B(g_input[19]), .Z(n19758) );
  XOR U19835 ( .A(n19857), .B(n19858), .Z(n19854) );
  AND U19836 ( .A(n19761), .B(n19859), .Z(n19858) );
  XNOR U19837 ( .A(n19728), .B(n19857), .Z(n19859) );
  XNOR U19838 ( .A(n19857), .B(g_input[18]), .Z(n19761) );
  XOR U19839 ( .A(n19860), .B(n19861), .Z(n19857) );
  AND U19840 ( .A(n19764), .B(n19862), .Z(n19861) );
  XNOR U19841 ( .A(n19728), .B(n19860), .Z(n19862) );
  XNOR U19842 ( .A(n19860), .B(g_input[17]), .Z(n19764) );
  XOR U19843 ( .A(n19863), .B(n19864), .Z(n19860) );
  AND U19844 ( .A(n19767), .B(n19865), .Z(n19864) );
  XNOR U19845 ( .A(n19728), .B(n19863), .Z(n19865) );
  XNOR U19846 ( .A(n19863), .B(g_input[16]), .Z(n19767) );
  XOR U19847 ( .A(n19866), .B(n19867), .Z(n19863) );
  AND U19848 ( .A(n19770), .B(n19868), .Z(n19867) );
  XNOR U19849 ( .A(n19728), .B(n19866), .Z(n19868) );
  XNOR U19850 ( .A(n19866), .B(g_input[15]), .Z(n19770) );
  XOR U19851 ( .A(n19869), .B(n19870), .Z(n19866) );
  AND U19852 ( .A(n19773), .B(n19871), .Z(n19870) );
  XNOR U19853 ( .A(n19728), .B(n19869), .Z(n19871) );
  XNOR U19854 ( .A(n19869), .B(g_input[14]), .Z(n19773) );
  XOR U19855 ( .A(n19872), .B(n19873), .Z(n19869) );
  AND U19856 ( .A(n19776), .B(n19874), .Z(n19873) );
  XNOR U19857 ( .A(n19728), .B(n19872), .Z(n19874) );
  XNOR U19858 ( .A(n19872), .B(g_input[13]), .Z(n19776) );
  XOR U19859 ( .A(n19875), .B(n19876), .Z(n19872) );
  AND U19860 ( .A(n19779), .B(n19877), .Z(n19876) );
  XNOR U19861 ( .A(n19728), .B(n19875), .Z(n19877) );
  XNOR U19862 ( .A(n19875), .B(g_input[12]), .Z(n19779) );
  XOR U19863 ( .A(n19878), .B(n19879), .Z(n19875) );
  AND U19864 ( .A(n19782), .B(n19880), .Z(n19879) );
  XNOR U19865 ( .A(n19728), .B(n19878), .Z(n19880) );
  XNOR U19866 ( .A(n19878), .B(g_input[11]), .Z(n19782) );
  XOR U19867 ( .A(n19881), .B(n19882), .Z(n19878) );
  AND U19868 ( .A(n19785), .B(n19883), .Z(n19882) );
  XNOR U19869 ( .A(n19728), .B(n19881), .Z(n19883) );
  XNOR U19870 ( .A(n19881), .B(g_input[10]), .Z(n19785) );
  XOR U19871 ( .A(n19884), .B(n19885), .Z(n19881) );
  AND U19872 ( .A(n19788), .B(n19886), .Z(n19885) );
  XNOR U19873 ( .A(n19728), .B(n19884), .Z(n19886) );
  XNOR U19874 ( .A(n19884), .B(g_input[9]), .Z(n19788) );
  XOR U19875 ( .A(n19887), .B(n19888), .Z(n19884) );
  AND U19876 ( .A(n19791), .B(n19889), .Z(n19888) );
  XNOR U19877 ( .A(n19728), .B(n19887), .Z(n19889) );
  XNOR U19878 ( .A(n19887), .B(g_input[8]), .Z(n19791) );
  XOR U19879 ( .A(n19890), .B(n19891), .Z(n19887) );
  AND U19880 ( .A(n19794), .B(n19892), .Z(n19891) );
  XNOR U19881 ( .A(n19728), .B(n19890), .Z(n19892) );
  IV U19882 ( .A(e_input[16]), .Z(n19728) );
  XNOR U19883 ( .A(n19890), .B(g_input[7]), .Z(n19794) );
  XOR U19884 ( .A(n19893), .B(n19894), .Z(n19890) );
  AND U19885 ( .A(n19797), .B(n19895), .Z(n19894) );
  XOR U19886 ( .A(e_input[15]), .B(n19893), .Z(n19895) );
  XNOR U19887 ( .A(n19893), .B(g_input[6]), .Z(n19797) );
  XOR U19888 ( .A(n19896), .B(n19897), .Z(n19893) );
  AND U19889 ( .A(n19800), .B(n19898), .Z(n19897) );
  XOR U19890 ( .A(e_input[14]), .B(n19896), .Z(n19898) );
  XNOR U19891 ( .A(n19896), .B(g_input[5]), .Z(n19800) );
  XOR U19892 ( .A(n19899), .B(n19900), .Z(n19896) );
  AND U19893 ( .A(n19803), .B(n19901), .Z(n19900) );
  XOR U19894 ( .A(e_input[13]), .B(n19899), .Z(n19901) );
  XNOR U19895 ( .A(n19899), .B(g_input[4]), .Z(n19803) );
  XOR U19896 ( .A(n19902), .B(n19903), .Z(n19899) );
  AND U19897 ( .A(n19806), .B(n19904), .Z(n19903) );
  XOR U19898 ( .A(e_input[12]), .B(n19902), .Z(n19904) );
  XNOR U19899 ( .A(n19902), .B(g_input[3]), .Z(n19806) );
  XOR U19900 ( .A(n19905), .B(n19906), .Z(n19902) );
  AND U19901 ( .A(n19809), .B(n19907), .Z(n19906) );
  XOR U19902 ( .A(e_input[11]), .B(n19905), .Z(n19907) );
  XNOR U19903 ( .A(n19905), .B(g_input[2]), .Z(n19809) );
  XNOR U19904 ( .A(n19908), .B(n19909), .Z(n19905) );
  NANDN U19905 ( .B(n19910), .A(n19911), .Z(n19908) );
  XOR U19906 ( .A(e_input[10]), .B(n19909), .Z(n19911) );
  XOR U19907 ( .A(n19813), .B(n19812), .Z(n19815) );
  XNOR U19908 ( .A(n19912), .B(n19811), .Z(n19812) );
  XOR U19909 ( .A(e_input[9]), .B(g_input[0]), .Z(n19811) );
  IV U19910 ( .A(n19912), .Z(n19813) );
  XOR U19911 ( .A(n19910), .B(e_input[10]), .Z(n19912) );
  XOR U19912 ( .A(n19909), .B(g_input[1]), .Z(n19910) );
  ANDN U19913 ( .A(e_input[9]), .B(g_input[0]), .Z(n19909) );
endmodule

