module AND(
	input A, B,
	output Z
);

endmodule

module NOR(
	input A, B,
	output Z
);

endmodule

module XOR(
	input A, B,
	output Z
);

endmodule

module XNOR(
	input A, B,
	output Z
);

endmodule

module IV(
	input A,
	output Z
);

endmodule

